magic
tech gf180mcuC
magscale 1 10
timestamp 1670119371
<< metal1 >>
rect 40450 56702 40462 56754
rect 40514 56751 40526 56754
rect 41010 56751 41022 56754
rect 40514 56705 41022 56751
rect 40514 56702 40526 56705
rect 41010 56702 41022 56705
rect 41074 56702 41086 56754
rect 37090 56590 37102 56642
rect 37154 56639 37166 56642
rect 37762 56639 37774 56642
rect 37154 56593 37774 56639
rect 37154 56590 37166 56593
rect 37762 56590 37774 56593
rect 37826 56590 37838 56642
rect 41122 56590 41134 56642
rect 41186 56639 41198 56642
rect 41682 56639 41694 56642
rect 41186 56593 41694 56639
rect 41186 56590 41198 56593
rect 41682 56590 41694 56593
rect 41746 56590 41758 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 4846 56306 4898 56318
rect 4846 56242 4898 56254
rect 9662 56306 9714 56318
rect 9662 56242 9714 56254
rect 11006 56306 11058 56318
rect 11006 56242 11058 56254
rect 13694 56306 13746 56318
rect 13694 56242 13746 56254
rect 14366 56306 14418 56318
rect 14366 56242 14418 56254
rect 16382 56306 16434 56318
rect 16382 56242 16434 56254
rect 19070 56306 19122 56318
rect 19070 56242 19122 56254
rect 19742 56306 19794 56318
rect 19742 56242 19794 56254
rect 21422 56306 21474 56318
rect 21422 56242 21474 56254
rect 22430 56306 22482 56318
rect 22430 56242 22482 56254
rect 27134 56306 27186 56318
rect 27134 56242 27186 56254
rect 28366 56306 28418 56318
rect 28366 56242 28418 56254
rect 29822 56306 29874 56318
rect 29822 56242 29874 56254
rect 31838 56306 31890 56318
rect 31838 56242 31890 56254
rect 33182 56306 33234 56318
rect 33182 56242 33234 56254
rect 33854 56306 33906 56318
rect 33854 56242 33906 56254
rect 37102 56306 37154 56318
rect 37102 56242 37154 56254
rect 37774 56306 37826 56318
rect 37774 56242 37826 56254
rect 38558 56306 38610 56318
rect 38558 56242 38610 56254
rect 39230 56306 39282 56318
rect 39230 56242 39282 56254
rect 41022 56306 41074 56318
rect 41022 56242 41074 56254
rect 41694 56306 41746 56318
rect 41694 56242 41746 56254
rect 43934 56306 43986 56318
rect 43934 56242 43986 56254
rect 45502 56306 45554 56318
rect 45502 56242 45554 56254
rect 47966 56306 48018 56318
rect 47966 56242 48018 56254
rect 48862 56306 48914 56318
rect 48862 56242 48914 56254
rect 49534 56306 49586 56318
rect 49534 56242 49586 56254
rect 1822 56194 1874 56206
rect 3042 56142 3054 56194
rect 3106 56142 3118 56194
rect 5842 56142 5854 56194
rect 5906 56142 5918 56194
rect 46050 56142 46062 56194
rect 46114 56142 46126 56194
rect 54898 56142 54910 56194
rect 54962 56142 54974 56194
rect 1822 56130 1874 56142
rect 15038 56082 15090 56094
rect 4162 56030 4174 56082
rect 4226 56030 4238 56082
rect 12786 56030 12798 56082
rect 12850 56030 12862 56082
rect 56802 56030 56814 56082
rect 56866 56030 56878 56082
rect 15038 56018 15090 56030
rect 54014 55970 54066 55982
rect 7186 55918 7198 55970
rect 7250 55918 7262 55970
rect 12002 55918 12014 55970
rect 12066 55918 12078 55970
rect 47170 55918 47182 55970
rect 47234 55918 47246 55970
rect 55906 55918 55918 55970
rect 55970 55918 55982 55970
rect 57362 55918 57374 55970
rect 57426 55918 57438 55970
rect 54014 55906 54066 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 5742 55410 5794 55422
rect 46274 55358 46286 55410
rect 46338 55358 46350 55410
rect 48402 55358 48414 55410
rect 48466 55358 48478 55410
rect 55122 55358 55134 55410
rect 55186 55358 55198 55410
rect 5742 55346 5794 55358
rect 3042 55246 3054 55298
rect 3106 55246 3118 55298
rect 45602 55246 45614 55298
rect 45666 55246 45678 55298
rect 3614 55186 3666 55198
rect 1922 55134 1934 55186
rect 1986 55134 1998 55186
rect 3614 55122 3666 55134
rect 4286 55186 4338 55198
rect 4286 55122 4338 55134
rect 13694 55186 13746 55198
rect 57374 55186 57426 55198
rect 56242 55134 56254 55186
rect 56306 55134 56318 55186
rect 13694 55122 13746 55134
rect 57374 55122 57426 55134
rect 57934 55186 57986 55198
rect 57934 55122 57986 55134
rect 4846 55074 4898 55086
rect 4846 55010 4898 55022
rect 48862 55074 48914 55086
rect 48862 55010 48914 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 2494 54738 2546 54750
rect 2494 54674 2546 54686
rect 3166 54738 3218 54750
rect 3166 54674 3218 54686
rect 56702 54738 56754 54750
rect 56702 54674 56754 54686
rect 58046 54738 58098 54750
rect 58046 54674 58098 54686
rect 1822 54626 1874 54638
rect 1822 54562 1874 54574
rect 52222 54626 52274 54638
rect 53554 54574 53566 54626
rect 53618 54574 53630 54626
rect 52222 54562 52274 54574
rect 51886 54514 51938 54526
rect 44482 54462 44494 54514
rect 44546 54462 44558 54514
rect 52882 54462 52894 54514
rect 52946 54462 52958 54514
rect 51886 54450 51938 54462
rect 3726 54402 3778 54414
rect 44942 54402 44994 54414
rect 56254 54402 56306 54414
rect 41570 54350 41582 54402
rect 41634 54350 41646 54402
rect 43698 54350 43710 54402
rect 43762 54350 43774 54402
rect 55682 54350 55694 54402
rect 55746 54350 55758 54402
rect 3726 54338 3778 54350
rect 44942 54338 44994 54350
rect 56254 54338 56306 54350
rect 55906 54238 55918 54290
rect 55970 54287 55982 54290
rect 56802 54287 56814 54290
rect 55970 54241 56814 54287
rect 55970 54238 55982 54241
rect 56802 54238 56814 54241
rect 56866 54238 56878 54290
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 43922 53790 43934 53842
rect 43986 53790 43998 53842
rect 50082 53790 50094 53842
rect 50146 53790 50158 53842
rect 44718 53730 44770 53742
rect 3042 53678 3054 53730
rect 3106 53678 3118 53730
rect 44146 53678 44158 53730
rect 44210 53678 44222 53730
rect 47282 53678 47294 53730
rect 47346 53678 47358 53730
rect 44718 53666 44770 53678
rect 50542 53618 50594 53630
rect 1922 53566 1934 53618
rect 1986 53566 1998 53618
rect 47954 53566 47966 53618
rect 48018 53566 48030 53618
rect 50542 53554 50594 53566
rect 3502 53506 3554 53518
rect 3502 53442 3554 53454
rect 46734 53506 46786 53518
rect 46734 53442 46786 53454
rect 58046 53506 58098 53518
rect 58046 53442 58098 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 44270 53170 44322 53182
rect 44270 53106 44322 53118
rect 44382 53170 44434 53182
rect 44382 53106 44434 53118
rect 45278 53170 45330 53182
rect 45278 53106 45330 53118
rect 1822 53058 1874 53070
rect 1822 52994 1874 53006
rect 45502 53058 45554 53070
rect 45502 52994 45554 53006
rect 48078 53058 48130 53070
rect 48078 52994 48130 53006
rect 58046 53058 58098 53070
rect 58046 52994 58098 53006
rect 44158 52946 44210 52958
rect 45614 52946 45666 52958
rect 44706 52894 44718 52946
rect 44770 52894 44782 52946
rect 44158 52882 44210 52894
rect 45614 52882 45666 52894
rect 48190 52946 48242 52958
rect 52994 52894 53006 52946
rect 53058 52894 53070 52946
rect 48190 52882 48242 52894
rect 48638 52834 48690 52846
rect 48638 52770 48690 52782
rect 49422 52834 49474 52846
rect 53454 52834 53506 52846
rect 50082 52782 50094 52834
rect 50146 52782 50158 52834
rect 52210 52782 52222 52834
rect 52274 52782 52286 52834
rect 49422 52770 49474 52782
rect 53454 52770 53506 52782
rect 48078 52722 48130 52734
rect 48402 52670 48414 52722
rect 48466 52719 48478 52722
rect 48626 52719 48638 52722
rect 48466 52673 48638 52719
rect 48466 52670 48478 52673
rect 48626 52670 48638 52673
rect 48690 52670 48702 52722
rect 48078 52658 48130 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 43262 52274 43314 52286
rect 39890 52222 39902 52274
rect 39954 52222 39966 52274
rect 45602 52222 45614 52274
rect 45666 52222 45678 52274
rect 53442 52222 53454 52274
rect 53506 52222 53518 52274
rect 55570 52222 55582 52274
rect 55634 52222 55646 52274
rect 43262 52210 43314 52222
rect 44830 52162 44882 52174
rect 48190 52162 48242 52174
rect 42018 52110 42030 52162
rect 42082 52110 42094 52162
rect 42802 52110 42814 52162
rect 42866 52110 42878 52162
rect 47954 52110 47966 52162
rect 48018 52110 48030 52162
rect 44830 52098 44882 52110
rect 48190 52098 48242 52110
rect 49086 52162 49138 52174
rect 56814 52162 56866 52174
rect 56242 52110 56254 52162
rect 56306 52110 56318 52162
rect 49086 52098 49138 52110
rect 56814 52098 56866 52110
rect 44494 52050 44546 52062
rect 44494 51986 44546 51998
rect 45950 52050 46002 52062
rect 45950 51986 46002 51998
rect 47294 52050 47346 52062
rect 47294 51986 47346 51998
rect 51326 52050 51378 52062
rect 51326 51986 51378 51998
rect 51662 52050 51714 52062
rect 51662 51986 51714 51998
rect 44046 51938 44098 51950
rect 44046 51874 44098 51886
rect 44606 51938 44658 51950
rect 44606 51874 44658 51886
rect 45502 51938 45554 51950
rect 45502 51874 45554 51886
rect 45726 51938 45778 51950
rect 45726 51874 45778 51886
rect 46398 51938 46450 51950
rect 46398 51874 46450 51886
rect 48750 51938 48802 51950
rect 48750 51874 48802 51886
rect 48974 51938 49026 51950
rect 48974 51874 49026 51886
rect 49646 51938 49698 51950
rect 49646 51874 49698 51886
rect 50094 51938 50146 51950
rect 50094 51874 50146 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 41918 51602 41970 51614
rect 41918 51538 41970 51550
rect 44494 51602 44546 51614
rect 44494 51538 44546 51550
rect 45614 51602 45666 51614
rect 45614 51538 45666 51550
rect 49422 51602 49474 51614
rect 49422 51538 49474 51550
rect 53454 51602 53506 51614
rect 53454 51538 53506 51550
rect 1822 51490 1874 51502
rect 1822 51426 1874 51438
rect 44046 51490 44098 51502
rect 44046 51426 44098 51438
rect 44718 51490 44770 51502
rect 44718 51426 44770 51438
rect 44830 51490 44882 51502
rect 44830 51426 44882 51438
rect 45838 51490 45890 51502
rect 45838 51426 45890 51438
rect 46622 51490 46674 51502
rect 46622 51426 46674 51438
rect 46734 51490 46786 51502
rect 46734 51426 46786 51438
rect 49646 51490 49698 51502
rect 49646 51426 49698 51438
rect 58046 51490 58098 51502
rect 58046 51426 58098 51438
rect 45950 51378 46002 51390
rect 41682 51326 41694 51378
rect 41746 51326 41758 51378
rect 45950 51314 46002 51326
rect 46398 51378 46450 51390
rect 49758 51378 49810 51390
rect 48066 51326 48078 51378
rect 48130 51326 48142 51378
rect 46398 51314 46450 51326
rect 49758 51314 49810 51326
rect 50206 51266 50258 51278
rect 48178 51214 48190 51266
rect 48242 51214 48254 51266
rect 50206 51202 50258 51214
rect 50654 51266 50706 51278
rect 50654 51202 50706 51214
rect 51326 51266 51378 51278
rect 51326 51202 51378 51214
rect 52558 51266 52610 51278
rect 52558 51202 52610 51214
rect 53006 51266 53058 51278
rect 53006 51202 53058 51214
rect 54798 51266 54850 51278
rect 54798 51202 54850 51214
rect 47618 51102 47630 51154
rect 47682 51102 47694 51154
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 49186 50766 49198 50818
rect 49250 50815 49262 50818
rect 49858 50815 49870 50818
rect 49250 50769 49870 50815
rect 49250 50766 49262 50769
rect 49858 50766 49870 50769
rect 49922 50766 49934 50818
rect 42926 50706 42978 50718
rect 49870 50706 49922 50718
rect 39554 50654 39566 50706
rect 39618 50654 39630 50706
rect 46274 50654 46286 50706
rect 46338 50654 46350 50706
rect 47618 50654 47630 50706
rect 47682 50654 47694 50706
rect 51762 50654 51774 50706
rect 51826 50654 51838 50706
rect 55122 50654 55134 50706
rect 55186 50654 55198 50706
rect 57250 50654 57262 50706
rect 57314 50654 57326 50706
rect 42926 50642 42978 50654
rect 49870 50642 49922 50654
rect 51438 50594 51490 50606
rect 42466 50542 42478 50594
rect 42530 50542 42542 50594
rect 46386 50542 46398 50594
rect 46450 50542 46462 50594
rect 47842 50542 47854 50594
rect 47906 50542 47918 50594
rect 52210 50542 52222 50594
rect 52274 50542 52286 50594
rect 57922 50542 57934 50594
rect 57986 50542 57998 50594
rect 51438 50530 51490 50542
rect 44718 50482 44770 50494
rect 41682 50430 41694 50482
rect 41746 50430 41758 50482
rect 44718 50418 44770 50430
rect 45502 50482 45554 50494
rect 45502 50418 45554 50430
rect 47182 50482 47234 50494
rect 47182 50418 47234 50430
rect 48974 50482 49026 50494
rect 48974 50418 49026 50430
rect 49422 50482 49474 50494
rect 49422 50418 49474 50430
rect 48638 50370 48690 50382
rect 48638 50306 48690 50318
rect 48862 50370 48914 50382
rect 48862 50306 48914 50318
rect 50318 50370 50370 50382
rect 50318 50306 50370 50318
rect 50878 50370 50930 50382
rect 50878 50306 50930 50318
rect 53342 50370 53394 50382
rect 53342 50306 53394 50318
rect 53790 50370 53842 50382
rect 53790 50306 53842 50318
rect 54350 50370 54402 50382
rect 54350 50306 54402 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 44494 50034 44546 50046
rect 44494 49970 44546 49982
rect 47294 50034 47346 50046
rect 47294 49970 47346 49982
rect 47406 50034 47458 50046
rect 47406 49970 47458 49982
rect 49422 50034 49474 50046
rect 49422 49970 49474 49982
rect 50430 50034 50482 50046
rect 50430 49970 50482 49982
rect 52110 50034 52162 50046
rect 52110 49970 52162 49982
rect 53454 50034 53506 50046
rect 53454 49970 53506 49982
rect 58046 50034 58098 50046
rect 58046 49970 58098 49982
rect 48638 49922 48690 49934
rect 48638 49858 48690 49870
rect 48750 49922 48802 49934
rect 48750 49858 48802 49870
rect 52894 49922 52946 49934
rect 52894 49858 52946 49870
rect 53006 49922 53058 49934
rect 53006 49858 53058 49870
rect 53678 49922 53730 49934
rect 53678 49858 53730 49870
rect 44382 49810 44434 49822
rect 44382 49746 44434 49758
rect 44606 49810 44658 49822
rect 44606 49746 44658 49758
rect 44942 49810 44994 49822
rect 44942 49746 44994 49758
rect 45614 49810 45666 49822
rect 47518 49810 47570 49822
rect 47966 49810 48018 49822
rect 45826 49758 45838 49810
rect 45890 49758 45902 49810
rect 47618 49758 47630 49810
rect 47682 49758 47694 49810
rect 45614 49746 45666 49758
rect 47518 49746 47570 49758
rect 47966 49746 48018 49758
rect 48414 49810 48466 49822
rect 48414 49746 48466 49758
rect 50990 49810 51042 49822
rect 51774 49810 51826 49822
rect 51538 49758 51550 49810
rect 51602 49758 51614 49810
rect 50990 49746 51042 49758
rect 51774 49746 51826 49758
rect 51998 49810 52050 49822
rect 51998 49746 52050 49758
rect 52670 49810 52722 49822
rect 52670 49746 52722 49758
rect 53790 49810 53842 49822
rect 56130 49758 56142 49810
rect 56194 49758 56206 49810
rect 53790 49746 53842 49758
rect 49870 49698 49922 49710
rect 49870 49634 49922 49646
rect 51886 49698 51938 49710
rect 51886 49634 51938 49646
rect 54238 49698 54290 49710
rect 56590 49698 56642 49710
rect 55346 49646 55358 49698
rect 55410 49646 55422 49698
rect 54238 49634 54290 49646
rect 56590 49634 56642 49646
rect 45502 49586 45554 49598
rect 49298 49534 49310 49586
rect 49362 49583 49374 49586
rect 50194 49583 50206 49586
rect 49362 49537 50206 49583
rect 49362 49534 49374 49537
rect 50194 49534 50206 49537
rect 50258 49534 50270 49586
rect 45502 49522 45554 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 47518 49250 47570 49262
rect 51102 49250 51154 49262
rect 48178 49198 48190 49250
rect 48242 49198 48254 49250
rect 47518 49186 47570 49198
rect 51102 49186 51154 49198
rect 53566 49250 53618 49262
rect 53566 49186 53618 49198
rect 42702 49138 42754 49150
rect 42702 49074 42754 49086
rect 48750 49138 48802 49150
rect 48750 49074 48802 49086
rect 49198 49138 49250 49150
rect 58034 49086 58046 49138
rect 58098 49086 58110 49138
rect 49198 49074 49250 49086
rect 43262 49026 43314 49038
rect 45838 49026 45890 49038
rect 41122 48974 41134 49026
rect 41186 48974 41198 49026
rect 44146 48974 44158 49026
rect 44210 48974 44222 49026
rect 44482 48974 44494 49026
rect 44546 48974 44558 49026
rect 43262 48962 43314 48974
rect 45838 48962 45890 48974
rect 46062 49026 46114 49038
rect 46062 48962 46114 48974
rect 48526 49026 48578 49038
rect 48526 48962 48578 48974
rect 50094 49026 50146 49038
rect 54574 49026 54626 49038
rect 50642 48974 50654 49026
rect 50706 48974 50718 49026
rect 51650 48974 51662 49026
rect 51714 48974 51726 49026
rect 52546 48974 52558 49026
rect 52610 48974 52622 49026
rect 55234 48974 55246 49026
rect 55298 48974 55310 49026
rect 50094 48962 50146 48974
rect 54574 48962 54626 48974
rect 41358 48914 41410 48926
rect 41358 48850 41410 48862
rect 44718 48914 44770 48926
rect 44718 48850 44770 48862
rect 45950 48914 46002 48926
rect 45950 48850 46002 48862
rect 46398 48914 46450 48926
rect 46398 48850 46450 48862
rect 46958 48914 47010 48926
rect 46958 48850 47010 48862
rect 47406 48914 47458 48926
rect 47406 48850 47458 48862
rect 50318 48914 50370 48926
rect 53678 48914 53730 48926
rect 50530 48862 50542 48914
rect 50594 48862 50606 48914
rect 52658 48862 52670 48914
rect 52722 48862 52734 48914
rect 55906 48862 55918 48914
rect 55970 48862 55982 48914
rect 50318 48850 50370 48862
rect 53678 48850 53730 48862
rect 42590 48802 42642 48814
rect 42590 48738 42642 48750
rect 42814 48802 42866 48814
rect 42814 48738 42866 48750
rect 47518 48802 47570 48814
rect 53566 48802 53618 48814
rect 51650 48750 51662 48802
rect 51714 48750 51726 48802
rect 47518 48738 47570 48750
rect 53566 48738 53618 48750
rect 54126 48802 54178 48814
rect 54126 48738 54178 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 49870 48466 49922 48478
rect 49870 48402 49922 48414
rect 50318 48466 50370 48478
rect 50318 48402 50370 48414
rect 52446 48466 52498 48478
rect 52446 48402 52498 48414
rect 52782 48466 52834 48478
rect 52782 48402 52834 48414
rect 57374 48466 57426 48478
rect 57374 48402 57426 48414
rect 41694 48354 41746 48366
rect 41694 48290 41746 48302
rect 47518 48354 47570 48366
rect 47518 48290 47570 48302
rect 48302 48354 48354 48366
rect 58046 48354 58098 48366
rect 53554 48302 53566 48354
rect 53618 48302 53630 48354
rect 53890 48302 53902 48354
rect 53954 48302 53966 48354
rect 55346 48302 55358 48354
rect 55410 48302 55422 48354
rect 48302 48290 48354 48302
rect 58046 48290 58098 48302
rect 42590 48242 42642 48254
rect 44718 48242 44770 48254
rect 46510 48242 46562 48254
rect 42354 48190 42366 48242
rect 42418 48190 42430 48242
rect 44258 48190 44270 48242
rect 44322 48190 44334 48242
rect 45826 48190 45838 48242
rect 45890 48190 45902 48242
rect 42590 48178 42642 48190
rect 44718 48178 44770 48190
rect 46510 48178 46562 48190
rect 46734 48242 46786 48254
rect 46734 48178 46786 48190
rect 47294 48242 47346 48254
rect 47294 48178 47346 48190
rect 51774 48242 51826 48254
rect 51774 48178 51826 48190
rect 51998 48242 52050 48254
rect 51998 48178 52050 48190
rect 53454 48242 53506 48254
rect 53454 48178 53506 48190
rect 54238 48242 54290 48254
rect 54238 48178 54290 48190
rect 44830 48130 44882 48142
rect 48750 48130 48802 48142
rect 47618 48078 47630 48130
rect 47682 48078 47694 48130
rect 44830 48066 44882 48078
rect 48750 48066 48802 48078
rect 49422 48130 49474 48142
rect 49422 48066 49474 48078
rect 50990 48130 51042 48142
rect 50990 48066 51042 48078
rect 51550 48130 51602 48142
rect 56354 48078 56366 48130
rect 56418 48078 56430 48130
rect 51550 48066 51602 48078
rect 48190 48018 48242 48030
rect 54462 48018 54514 48030
rect 49410 47966 49422 48018
rect 49474 48015 49486 48018
rect 50194 48015 50206 48018
rect 49474 47969 50206 48015
rect 49474 47966 49486 47969
rect 50194 47966 50206 47969
rect 50258 47966 50270 48018
rect 48190 47954 48242 47966
rect 54462 47954 54514 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 44270 47682 44322 47694
rect 42578 47630 42590 47682
rect 42642 47630 42654 47682
rect 44270 47618 44322 47630
rect 51998 47682 52050 47694
rect 51998 47618 52050 47630
rect 45502 47570 45554 47582
rect 49310 47570 49362 47582
rect 43138 47518 43150 47570
rect 43202 47518 43214 47570
rect 46386 47518 46398 47570
rect 46450 47518 46462 47570
rect 45502 47506 45554 47518
rect 49310 47506 49362 47518
rect 49758 47570 49810 47582
rect 49758 47506 49810 47518
rect 50654 47570 50706 47582
rect 50654 47506 50706 47518
rect 51102 47570 51154 47582
rect 51102 47506 51154 47518
rect 53342 47570 53394 47582
rect 54450 47518 54462 47570
rect 54514 47518 54526 47570
rect 55122 47518 55134 47570
rect 55186 47518 55198 47570
rect 57250 47518 57262 47570
rect 57314 47518 57326 47570
rect 53342 47506 53394 47518
rect 44382 47458 44434 47470
rect 47406 47458 47458 47470
rect 43362 47406 43374 47458
rect 43426 47406 43438 47458
rect 46162 47406 46174 47458
rect 46226 47406 46238 47458
rect 44382 47394 44434 47406
rect 47406 47394 47458 47406
rect 48078 47458 48130 47470
rect 48078 47394 48130 47406
rect 51774 47458 51826 47470
rect 54126 47458 54178 47470
rect 53890 47406 53902 47458
rect 53954 47406 53966 47458
rect 51774 47394 51826 47406
rect 54126 47394 54178 47406
rect 54350 47458 54402 47470
rect 57922 47406 57934 47458
rect 57986 47406 57998 47458
rect 54350 47394 54402 47406
rect 47854 47346 47906 47358
rect 47854 47282 47906 47294
rect 48862 47346 48914 47358
rect 48862 47282 48914 47294
rect 54462 47346 54514 47358
rect 54462 47282 54514 47294
rect 1822 47234 1874 47246
rect 1822 47170 1874 47182
rect 44270 47234 44322 47246
rect 44270 47170 44322 47182
rect 46958 47234 47010 47246
rect 46958 47170 47010 47182
rect 47630 47234 47682 47246
rect 47630 47170 47682 47182
rect 48526 47234 48578 47246
rect 48526 47170 48578 47182
rect 48750 47234 48802 47246
rect 48750 47170 48802 47182
rect 50206 47234 50258 47246
rect 52322 47182 52334 47234
rect 52386 47182 52398 47234
rect 50206 47170 50258 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 46958 46898 47010 46910
rect 46958 46834 47010 46846
rect 48190 46898 48242 46910
rect 48190 46834 48242 46846
rect 48302 46898 48354 46910
rect 48302 46834 48354 46846
rect 51214 46898 51266 46910
rect 51214 46834 51266 46846
rect 51438 46898 51490 46910
rect 51438 46834 51490 46846
rect 51550 46898 51602 46910
rect 51550 46834 51602 46846
rect 53678 46898 53730 46910
rect 53678 46834 53730 46846
rect 54798 46898 54850 46910
rect 54798 46834 54850 46846
rect 55806 46898 55858 46910
rect 55806 46834 55858 46846
rect 56254 46898 56306 46910
rect 56254 46834 56306 46846
rect 57486 46898 57538 46910
rect 57486 46834 57538 46846
rect 46174 46786 46226 46798
rect 46174 46722 46226 46734
rect 47070 46786 47122 46798
rect 47070 46722 47122 46734
rect 52334 46786 52386 46798
rect 52334 46722 52386 46734
rect 53006 46786 53058 46798
rect 53006 46722 53058 46734
rect 53118 46786 53170 46798
rect 53118 46722 53170 46734
rect 54574 46786 54626 46798
rect 54574 46722 54626 46734
rect 58046 46786 58098 46798
rect 58046 46722 58098 46734
rect 46510 46674 46562 46686
rect 48526 46674 48578 46686
rect 49982 46674 50034 46686
rect 47282 46622 47294 46674
rect 47346 46622 47358 46674
rect 47506 46622 47518 46674
rect 47570 46622 47582 46674
rect 48738 46622 48750 46674
rect 48802 46622 48814 46674
rect 46510 46610 46562 46622
rect 48526 46610 48578 46622
rect 49982 46610 50034 46622
rect 50206 46674 50258 46686
rect 52222 46674 52274 46686
rect 50978 46622 50990 46674
rect 51042 46622 51054 46674
rect 50206 46610 50258 46622
rect 52222 46610 52274 46622
rect 52558 46674 52610 46686
rect 52558 46610 52610 46622
rect 53342 46674 53394 46686
rect 53342 46610 53394 46622
rect 55470 46674 55522 46686
rect 55470 46610 55522 46622
rect 48414 46562 48466 46574
rect 48414 46498 48466 46510
rect 51326 46562 51378 46574
rect 51326 46498 51378 46510
rect 56702 46562 56754 46574
rect 56702 46498 56754 46510
rect 54910 46450 54962 46462
rect 49634 46398 49646 46450
rect 49698 46398 49710 46450
rect 56018 46398 56030 46450
rect 56082 46447 56094 46450
rect 56690 46447 56702 46450
rect 56082 46401 56702 46447
rect 56082 46398 56094 46401
rect 56690 46398 56702 46401
rect 56754 46398 56766 46450
rect 54910 46386 54962 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 50990 46114 51042 46126
rect 55010 46062 55022 46114
rect 55074 46111 55086 46114
rect 56018 46111 56030 46114
rect 55074 46065 56030 46111
rect 55074 46062 55086 46065
rect 56018 46062 56030 46065
rect 56082 46062 56094 46114
rect 50990 46050 51042 46062
rect 42926 46002 42978 46014
rect 42926 45938 42978 45950
rect 47182 46002 47234 46014
rect 47182 45938 47234 45950
rect 50094 46002 50146 46014
rect 50094 45938 50146 45950
rect 50766 46002 50818 46014
rect 50766 45938 50818 45950
rect 51998 46002 52050 46014
rect 51998 45938 52050 45950
rect 54462 46002 54514 46014
rect 54462 45938 54514 45950
rect 54910 46002 54962 46014
rect 54910 45938 54962 45950
rect 55918 46002 55970 46014
rect 55918 45938 55970 45950
rect 57374 46002 57426 46014
rect 57374 45938 57426 45950
rect 47294 45890 47346 45902
rect 48750 45890 48802 45902
rect 48178 45838 48190 45890
rect 48242 45838 48254 45890
rect 47294 45826 47346 45838
rect 48750 45826 48802 45838
rect 51886 45890 51938 45902
rect 51886 45826 51938 45838
rect 52110 45890 52162 45902
rect 52110 45826 52162 45838
rect 52334 45890 52386 45902
rect 52334 45826 52386 45838
rect 53454 45890 53506 45902
rect 53454 45826 53506 45838
rect 53678 45890 53730 45902
rect 53678 45826 53730 45838
rect 42814 45778 42866 45790
rect 42814 45714 42866 45726
rect 43150 45778 43202 45790
rect 43150 45714 43202 45726
rect 43374 45778 43426 45790
rect 43374 45714 43426 45726
rect 46174 45778 46226 45790
rect 46174 45714 46226 45726
rect 48414 45778 48466 45790
rect 54014 45778 54066 45790
rect 48626 45726 48638 45778
rect 48690 45726 48702 45778
rect 48414 45714 48466 45726
rect 54014 45714 54066 45726
rect 1822 45666 1874 45678
rect 1822 45602 1874 45614
rect 2494 45666 2546 45678
rect 2494 45602 2546 45614
rect 46286 45666 46338 45678
rect 46286 45602 46338 45614
rect 47742 45666 47794 45678
rect 47742 45602 47794 45614
rect 49198 45666 49250 45678
rect 49198 45602 49250 45614
rect 49646 45666 49698 45678
rect 53678 45666 53730 45678
rect 51314 45614 51326 45666
rect 51378 45614 51390 45666
rect 49646 45602 49698 45614
rect 53678 45602 53730 45614
rect 55582 45666 55634 45678
rect 55582 45602 55634 45614
rect 58046 45666 58098 45678
rect 58046 45602 58098 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 46286 45330 46338 45342
rect 46286 45266 46338 45278
rect 46398 45330 46450 45342
rect 46398 45266 46450 45278
rect 49534 45330 49586 45342
rect 49534 45266 49586 45278
rect 50766 45330 50818 45342
rect 50766 45266 50818 45278
rect 1822 45218 1874 45230
rect 1822 45154 1874 45166
rect 43598 45218 43650 45230
rect 55246 45218 55298 45230
rect 48290 45166 48302 45218
rect 48354 45166 48366 45218
rect 43598 45154 43650 45166
rect 55246 45154 55298 45166
rect 58046 45218 58098 45230
rect 58046 45154 58098 45166
rect 43710 45106 43762 45118
rect 46510 45106 46562 45118
rect 55806 45106 55858 45118
rect 42690 45054 42702 45106
rect 42754 45054 42766 45106
rect 44258 45054 44270 45106
rect 44322 45054 44334 45106
rect 47730 45054 47742 45106
rect 47794 45054 47806 45106
rect 48178 45054 48190 45106
rect 48242 45054 48254 45106
rect 51874 45054 51886 45106
rect 51938 45054 51950 45106
rect 53442 45054 53454 45106
rect 53506 45054 53518 45106
rect 54450 45054 54462 45106
rect 54514 45054 54526 45106
rect 43710 45042 43762 45054
rect 46510 45042 46562 45054
rect 55806 45042 55858 45054
rect 56366 45106 56418 45118
rect 56366 45042 56418 45054
rect 42030 44994 42082 45006
rect 45054 44994 45106 45006
rect 42802 44942 42814 44994
rect 42866 44942 42878 44994
rect 42030 44930 42082 44942
rect 45054 44930 45106 44942
rect 46062 44994 46114 45006
rect 52334 44994 52386 45006
rect 48514 44942 48526 44994
rect 48578 44942 48590 44994
rect 51986 44942 51998 44994
rect 52050 44942 52062 44994
rect 53330 44942 53342 44994
rect 53394 44942 53406 44994
rect 46062 44930 46114 44942
rect 52334 44930 52386 44942
rect 45614 44882 45666 44894
rect 45614 44818 45666 44830
rect 45838 44882 45890 44894
rect 45838 44818 45890 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 43374 44546 43426 44558
rect 43374 44482 43426 44494
rect 43710 44546 43762 44558
rect 43710 44482 43762 44494
rect 44718 44546 44770 44558
rect 48178 44494 48190 44546
rect 48242 44494 48254 44546
rect 44718 44482 44770 44494
rect 45502 44434 45554 44446
rect 45502 44370 45554 44382
rect 47070 44434 47122 44446
rect 47070 44370 47122 44382
rect 51438 44434 51490 44446
rect 55010 44382 55022 44434
rect 55074 44382 55086 44434
rect 51438 44370 51490 44382
rect 44606 44322 44658 44334
rect 44606 44258 44658 44270
rect 45614 44322 45666 44334
rect 49310 44322 49362 44334
rect 52782 44322 52834 44334
rect 45938 44270 45950 44322
rect 46002 44270 46014 44322
rect 48626 44270 48638 44322
rect 48690 44270 48702 44322
rect 49634 44270 49646 44322
rect 49698 44270 49710 44322
rect 52434 44270 52446 44322
rect 52498 44270 52510 44322
rect 45614 44258 45666 44270
rect 49310 44258 49362 44270
rect 52782 44258 52834 44270
rect 53342 44322 53394 44334
rect 53342 44258 53394 44270
rect 53902 44322 53954 44334
rect 57922 44270 57934 44322
rect 57986 44270 57998 44322
rect 53902 44258 53954 44270
rect 43486 44210 43538 44222
rect 43486 44146 43538 44158
rect 44494 44210 44546 44222
rect 52222 44210 52274 44222
rect 48402 44158 48414 44210
rect 48466 44158 48478 44210
rect 44494 44146 44546 44158
rect 52222 44146 52274 44158
rect 52670 44210 52722 44222
rect 52670 44146 52722 44158
rect 53790 44210 53842 44222
rect 57250 44158 57262 44210
rect 57314 44158 57326 44210
rect 53790 44146 53842 44158
rect 53566 44098 53618 44110
rect 53566 44034 53618 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 44046 43762 44098 43774
rect 44046 43698 44098 43710
rect 52334 43762 52386 43774
rect 52334 43698 52386 43710
rect 45502 43650 45554 43662
rect 45502 43586 45554 43598
rect 48750 43650 48802 43662
rect 48750 43586 48802 43598
rect 52558 43650 52610 43662
rect 52558 43586 52610 43598
rect 53566 43650 53618 43662
rect 53566 43586 53618 43598
rect 57598 43650 57650 43662
rect 57598 43586 57650 43598
rect 48526 43538 48578 43550
rect 45714 43486 45726 43538
rect 45778 43486 45790 43538
rect 46162 43486 46174 43538
rect 46226 43486 46238 43538
rect 47842 43486 47854 43538
rect 47906 43486 47918 43538
rect 48526 43474 48578 43486
rect 52670 43538 52722 43550
rect 52670 43474 52722 43486
rect 53118 43538 53170 43550
rect 53118 43474 53170 43486
rect 50430 43426 50482 43438
rect 50430 43362 50482 43374
rect 50878 43426 50930 43438
rect 50878 43362 50930 43374
rect 51326 43426 51378 43438
rect 51326 43362 51378 43374
rect 51774 43426 51826 43438
rect 51774 43362 51826 43374
rect 58046 43426 58098 43438
rect 58046 43362 58098 43374
rect 52882 43262 52894 43314
rect 52946 43311 52958 43314
rect 53442 43311 53454 43314
rect 52946 43265 53454 43311
rect 52946 43262 52958 43265
rect 53442 43262 53454 43265
rect 53506 43262 53518 43314
rect 57250 43262 57262 43314
rect 57314 43311 57326 43314
rect 58034 43311 58046 43314
rect 57314 43265 58046 43311
rect 57314 43262 57326 43265
rect 58034 43262 58046 43265
rect 58098 43262 58110 43314
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 53454 42978 53506 42990
rect 50194 42926 50206 42978
rect 50258 42975 50270 42978
rect 50978 42975 50990 42978
rect 50258 42929 50990 42975
rect 50258 42926 50270 42929
rect 50978 42926 50990 42929
rect 51042 42926 51054 42978
rect 53454 42914 53506 42926
rect 46286 42866 46338 42878
rect 43026 42814 43038 42866
rect 43090 42814 43102 42866
rect 46286 42802 46338 42814
rect 48526 42866 48578 42878
rect 50878 42866 50930 42878
rect 49410 42814 49422 42866
rect 49474 42814 49486 42866
rect 56354 42814 56366 42866
rect 56418 42814 56430 42866
rect 48526 42802 48578 42814
rect 50878 42802 50930 42814
rect 43598 42754 43650 42766
rect 40114 42702 40126 42754
rect 40178 42702 40190 42754
rect 43598 42690 43650 42702
rect 48750 42754 48802 42766
rect 49534 42754 49586 42766
rect 49298 42702 49310 42754
rect 49362 42702 49374 42754
rect 48750 42690 48802 42702
rect 49534 42690 49586 42702
rect 49982 42642 50034 42654
rect 40786 42590 40798 42642
rect 40850 42590 40862 42642
rect 48962 42590 48974 42642
rect 49026 42639 49038 42642
rect 49186 42639 49198 42642
rect 49026 42593 49198 42639
rect 49026 42590 49038 42593
rect 49186 42590 49198 42593
rect 49250 42590 49262 42642
rect 49982 42578 50034 42590
rect 51550 42642 51602 42654
rect 51550 42578 51602 42590
rect 52222 42642 52274 42654
rect 52222 42578 52274 42590
rect 53678 42642 53730 42654
rect 53678 42578 53730 42590
rect 54238 42642 54290 42654
rect 55234 42590 55246 42642
rect 55298 42590 55310 42642
rect 54238 42578 54290 42590
rect 39454 42530 39506 42542
rect 39454 42466 39506 42478
rect 46174 42530 46226 42542
rect 46174 42466 46226 42478
rect 46398 42530 46450 42542
rect 46398 42466 46450 42478
rect 46622 42530 46674 42542
rect 46622 42466 46674 42478
rect 48078 42530 48130 42542
rect 48078 42466 48130 42478
rect 48190 42530 48242 42542
rect 48190 42466 48242 42478
rect 48302 42530 48354 42542
rect 48302 42466 48354 42478
rect 49758 42530 49810 42542
rect 49758 42466 49810 42478
rect 50430 42530 50482 42542
rect 50430 42466 50482 42478
rect 51662 42530 51714 42542
rect 51662 42466 51714 42478
rect 52334 42530 52386 42542
rect 52334 42466 52386 42478
rect 53566 42530 53618 42542
rect 53566 42466 53618 42478
rect 56814 42530 56866 42542
rect 56814 42466 56866 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 52770 42142 52782 42194
rect 52834 42142 52846 42194
rect 47742 42082 47794 42094
rect 47742 42018 47794 42030
rect 49646 42082 49698 42094
rect 49646 42018 49698 42030
rect 49870 42082 49922 42094
rect 54238 42082 54290 42094
rect 51202 42030 51214 42082
rect 51266 42030 51278 42082
rect 49870 42018 49922 42030
rect 54238 42018 54290 42030
rect 46734 41970 46786 41982
rect 53678 41970 53730 41982
rect 46386 41918 46398 41970
rect 46450 41918 46462 41970
rect 48402 41918 48414 41970
rect 48466 41918 48478 41970
rect 52434 41918 52446 41970
rect 52498 41918 52510 41970
rect 46734 41906 46786 41918
rect 53678 41906 53730 41918
rect 54350 41970 54402 41982
rect 54350 41906 54402 41918
rect 46846 41858 46898 41870
rect 50318 41858 50370 41870
rect 53902 41858 53954 41870
rect 48626 41806 48638 41858
rect 48690 41806 48702 41858
rect 49522 41806 49534 41858
rect 49586 41806 49598 41858
rect 50978 41806 50990 41858
rect 51042 41806 51054 41858
rect 46846 41794 46898 41806
rect 50318 41794 50370 41806
rect 53902 41794 53954 41806
rect 54126 41858 54178 41870
rect 54126 41794 54178 41806
rect 54574 41746 54626 41758
rect 54574 41682 54626 41694
rect 54798 41746 54850 41758
rect 54798 41682 54850 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 47406 41410 47458 41422
rect 47406 41346 47458 41358
rect 49086 41410 49138 41422
rect 49086 41346 49138 41358
rect 49646 41410 49698 41422
rect 49646 41346 49698 41358
rect 50990 41410 51042 41422
rect 50990 41346 51042 41358
rect 52334 41410 52386 41422
rect 52658 41358 52670 41410
rect 52722 41358 52734 41410
rect 52334 41346 52386 41358
rect 45726 41298 45778 41310
rect 45726 41234 45778 41246
rect 50206 41298 50258 41310
rect 50206 41234 50258 41246
rect 51550 41298 51602 41310
rect 51550 41234 51602 41246
rect 52110 41298 52162 41310
rect 52110 41234 52162 41246
rect 53454 41298 53506 41310
rect 53454 41234 53506 41246
rect 53902 41298 53954 41310
rect 53902 41234 53954 41246
rect 54686 41298 54738 41310
rect 55122 41246 55134 41298
rect 55186 41246 55198 41298
rect 57250 41246 57262 41298
rect 57314 41246 57326 41298
rect 54686 41234 54738 41246
rect 46622 41186 46674 41198
rect 46386 41134 46398 41186
rect 46450 41134 46462 41186
rect 46622 41122 46674 41134
rect 47294 41186 47346 41198
rect 47294 41122 47346 41134
rect 48078 41186 48130 41198
rect 48078 41122 48130 41134
rect 48302 41186 48354 41198
rect 48302 41122 48354 41134
rect 48414 41186 48466 41198
rect 48414 41122 48466 41134
rect 48862 41186 48914 41198
rect 48862 41122 48914 41134
rect 49758 41186 49810 41198
rect 49758 41122 49810 41134
rect 51102 41186 51154 41198
rect 57922 41134 57934 41186
rect 57986 41134 57998 41186
rect 51102 41122 51154 41134
rect 47406 41074 47458 41086
rect 47406 41010 47458 41022
rect 49646 41074 49698 41086
rect 49646 41010 49698 41022
rect 50990 41074 51042 41086
rect 50990 41010 51042 41022
rect 1822 40962 1874 40974
rect 1822 40898 1874 40910
rect 2494 40962 2546 40974
rect 2494 40898 2546 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 44942 40626 44994 40638
rect 44942 40562 44994 40574
rect 46286 40626 46338 40638
rect 46286 40562 46338 40574
rect 46734 40626 46786 40638
rect 46734 40562 46786 40574
rect 48302 40626 48354 40638
rect 48302 40562 48354 40574
rect 48638 40626 48690 40638
rect 48638 40562 48690 40574
rect 50766 40626 50818 40638
rect 50766 40562 50818 40574
rect 51326 40626 51378 40638
rect 51326 40562 51378 40574
rect 51662 40626 51714 40638
rect 51662 40562 51714 40574
rect 52222 40626 52274 40638
rect 52222 40562 52274 40574
rect 1822 40514 1874 40526
rect 1822 40450 1874 40462
rect 46958 40514 47010 40526
rect 46958 40450 47010 40462
rect 47070 40514 47122 40526
rect 47070 40450 47122 40462
rect 47966 40514 48018 40526
rect 47966 40450 48018 40462
rect 48078 40514 48130 40526
rect 48078 40450 48130 40462
rect 49646 40514 49698 40526
rect 49646 40450 49698 40462
rect 49758 40514 49810 40526
rect 58046 40514 58098 40526
rect 56018 40462 56030 40514
rect 56082 40462 56094 40514
rect 49758 40450 49810 40462
rect 58046 40450 58098 40462
rect 40910 40402 40962 40414
rect 49982 40402 50034 40414
rect 41682 40350 41694 40402
rect 41746 40350 41758 40402
rect 42354 40350 42366 40402
rect 42418 40350 42430 40402
rect 40910 40338 40962 40350
rect 49982 40338 50034 40350
rect 50318 40402 50370 40414
rect 55122 40350 55134 40402
rect 55186 40350 55198 40402
rect 50318 40338 50370 40350
rect 44482 40238 44494 40290
rect 44546 40238 44558 40290
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 47406 39730 47458 39742
rect 47406 39666 47458 39678
rect 48414 39730 48466 39742
rect 50878 39730 50930 39742
rect 50306 39678 50318 39730
rect 50370 39678 50382 39730
rect 48414 39666 48466 39678
rect 50878 39666 50930 39678
rect 49970 39566 49982 39618
rect 50034 39566 50046 39618
rect 49422 39506 49474 39518
rect 49422 39442 49474 39454
rect 1822 39394 1874 39406
rect 1822 39330 1874 39342
rect 58046 39394 58098 39406
rect 58046 39330 58098 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 49534 38946 49586 38958
rect 49534 38882 49586 38894
rect 49746 38782 49758 38834
rect 49810 38782 49822 38834
rect 53666 38782 53678 38834
rect 53730 38782 53742 38834
rect 54238 38722 54290 38734
rect 50754 38670 50766 38722
rect 50818 38670 50830 38722
rect 52882 38670 52894 38722
rect 52946 38670 52958 38722
rect 54238 38658 54290 38670
rect 54574 38722 54626 38734
rect 54574 38658 54626 38670
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 53442 38110 53454 38162
rect 53506 38110 53518 38162
rect 56354 37998 56366 38050
rect 56418 37998 56430 38050
rect 55570 37886 55582 37938
rect 55634 37886 55646 37938
rect 56814 37826 56866 37838
rect 56814 37762 56866 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 53566 37490 53618 37502
rect 53566 37426 53618 37438
rect 54014 37378 54066 37390
rect 54014 37314 54066 37326
rect 54350 37378 54402 37390
rect 56242 37326 56254 37378
rect 56306 37326 56318 37378
rect 54350 37314 54402 37326
rect 57374 37154 57426 37166
rect 55122 37102 55134 37154
rect 55186 37102 55198 37154
rect 57374 37090 57426 37102
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 48290 36542 48302 36594
rect 48354 36542 48366 36594
rect 50418 36542 50430 36594
rect 50482 36542 50494 36594
rect 50878 36482 50930 36494
rect 47506 36430 47518 36482
rect 47570 36430 47582 36482
rect 50878 36418 50930 36430
rect 54898 36318 54910 36370
rect 54962 36318 54974 36370
rect 55246 36258 55298 36270
rect 55246 36194 55298 36206
rect 55806 36258 55858 36270
rect 55806 36194 55858 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 1822 35810 1874 35822
rect 1822 35746 1874 35758
rect 56130 35646 56142 35698
rect 56194 35646 56206 35698
rect 55346 35534 55358 35586
rect 55410 35534 55422 35586
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 54574 35026 54626 35038
rect 55906 34974 55918 35026
rect 55970 34974 55982 35026
rect 58034 34974 58046 35026
rect 58098 34974 58110 35026
rect 54574 34962 54626 34974
rect 55122 34862 55134 34914
rect 55186 34862 55198 34914
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 1822 31554 1874 31566
rect 1822 31490 1874 31502
rect 2494 31554 2546 31566
rect 2494 31490 2546 31502
rect 57374 31554 57426 31566
rect 57374 31490 57426 31502
rect 58046 31554 58098 31566
rect 58046 31490 58098 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 58046 31106 58098 31118
rect 58046 31042 58098 31054
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 1822 28418 1874 28430
rect 1822 28354 1874 28366
rect 58046 28418 58098 28430
rect 58046 28354 58098 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 1822 26850 1874 26862
rect 1822 26786 1874 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 42814 26514 42866 26526
rect 42814 26450 42866 26462
rect 42254 26402 42306 26414
rect 42254 26338 42306 26350
rect 42018 26238 42030 26290
rect 42082 26238 42094 26290
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 43934 25618 43986 25630
rect 40450 25566 40462 25618
rect 40514 25566 40526 25618
rect 42578 25566 42590 25618
rect 42642 25566 42654 25618
rect 43934 25554 43986 25566
rect 3042 25454 3054 25506
rect 3106 25454 3118 25506
rect 43362 25454 43374 25506
rect 43426 25454 43438 25506
rect 1922 25342 1934 25394
rect 1986 25342 1998 25394
rect 3614 25282 3666 25294
rect 3614 25218 3666 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 58046 24834 58098 24846
rect 58046 24770 58098 24782
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 1822 23266 1874 23278
rect 56242 23214 56254 23266
rect 56306 23214 56318 23266
rect 1822 23202 1874 23214
rect 57374 23042 57426 23054
rect 55122 22990 55134 23042
rect 55186 22990 55198 23042
rect 57374 22978 57426 22990
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 1822 22146 1874 22158
rect 1822 22082 1874 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 1822 21698 1874 21710
rect 1822 21634 1874 21646
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 1822 20130 1874 20142
rect 56242 20078 56254 20130
rect 56306 20078 56318 20130
rect 1822 20066 1874 20078
rect 57374 19906 57426 19918
rect 54898 19854 54910 19906
rect 54962 19854 54974 19906
rect 57374 19842 57426 19854
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 1822 18562 1874 18574
rect 1822 18498 1874 18510
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 1822 16994 1874 17006
rect 1822 16930 1874 16942
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 58046 15874 58098 15886
rect 58046 15810 58098 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 1822 15426 1874 15438
rect 1822 15362 1874 15374
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 1822 14306 1874 14318
rect 1822 14242 1874 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 58046 13858 58098 13870
rect 58046 13794 58098 13806
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 1822 12738 1874 12750
rect 1822 12674 1874 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 58046 11170 58098 11182
rect 58046 11106 58098 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 1822 10722 1874 10734
rect 1822 10658 1874 10670
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 1822 9602 1874 9614
rect 1822 9538 1874 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 1822 6466 1874 6478
rect 1822 6402 1874 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 58046 6018 58098 6030
rect 58046 5954 58098 5966
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 1822 4898 1874 4910
rect 1822 4834 1874 4846
rect 58046 4898 58098 4910
rect 58046 4834 58098 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 50766 4562 50818 4574
rect 50766 4498 50818 4510
rect 1822 4450 1874 4462
rect 1822 4386 1874 4398
rect 12350 4450 12402 4462
rect 58046 4450 58098 4462
rect 56242 4398 56254 4450
rect 56306 4398 56318 4450
rect 12350 4386 12402 4398
rect 58046 4386 58098 4398
rect 13022 4226 13074 4238
rect 57374 4226 57426 4238
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 13022 4162 13074 4174
rect 57374 4162 57426 4174
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 12786 3614 12798 3666
rect 12850 3614 12862 3666
rect 30706 3614 30718 3666
rect 30770 3614 30782 3666
rect 50530 3502 50542 3554
rect 50594 3502 50606 3554
rect 28590 3442 28642 3454
rect 11554 3390 11566 3442
rect 11618 3390 11630 3442
rect 29362 3390 29374 3442
rect 29426 3390 29438 3442
rect 49410 3390 49422 3442
rect 49474 3390 49486 3442
rect 28590 3378 28642 3390
rect 1822 3330 1874 3342
rect 1822 3266 1874 3278
rect 2494 3330 2546 3342
rect 2494 3266 2546 3278
rect 3614 3330 3666 3342
rect 3614 3266 3666 3278
rect 4286 3330 4338 3342
rect 4286 3266 4338 3278
rect 13582 3330 13634 3342
rect 13582 3266 13634 3278
rect 15038 3330 15090 3342
rect 15038 3266 15090 3278
rect 16382 3330 16434 3342
rect 16382 3266 16434 3278
rect 19070 3330 19122 3342
rect 19070 3266 19122 3278
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 23102 3330 23154 3342
rect 23102 3266 23154 3278
rect 24446 3330 24498 3342
rect 24446 3266 24498 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 37102 3330 37154 3342
rect 37102 3266 37154 3278
rect 39230 3330 39282 3342
rect 39230 3266 39282 3278
rect 39902 3330 39954 3342
rect 39902 3266 39954 3278
rect 46622 3330 46674 3342
rect 46622 3266 46674 3278
rect 47294 3330 47346 3342
rect 47294 3266 47346 3278
rect 48078 3330 48130 3342
rect 48078 3266 48130 3278
rect 51102 3330 51154 3342
rect 51102 3266 51154 3278
rect 51774 3330 51826 3342
rect 51774 3266 51826 3278
rect 55918 3330 55970 3342
rect 55918 3266 55970 3278
rect 56702 3330 56754 3342
rect 56702 3266 56754 3278
rect 57934 3330 57986 3342
rect 57934 3266 57986 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
rect 32386 1710 32398 1762
rect 32450 1759 32462 1762
rect 33170 1759 33182 1762
rect 32450 1713 33182 1759
rect 32450 1710 32462 1713
rect 33170 1710 33182 1713
rect 33234 1710 33246 1762
rect 50530 1710 50542 1762
rect 50594 1759 50606 1762
rect 51090 1759 51102 1762
rect 50594 1713 51102 1759
rect 50594 1710 50606 1713
rect 51090 1710 51102 1713
rect 51154 1710 51166 1762
rect 55906 1710 55918 1762
rect 55970 1759 55982 1762
rect 56690 1759 56702 1762
rect 55970 1713 56702 1759
rect 55970 1710 55982 1713
rect 56690 1710 56702 1713
rect 56754 1710 56766 1762
<< via1 >>
rect 40462 56702 40514 56754
rect 41022 56702 41074 56754
rect 37102 56590 37154 56642
rect 37774 56590 37826 56642
rect 41134 56590 41186 56642
rect 41694 56590 41746 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4846 56254 4898 56306
rect 9662 56254 9714 56306
rect 11006 56254 11058 56306
rect 13694 56254 13746 56306
rect 14366 56254 14418 56306
rect 16382 56254 16434 56306
rect 19070 56254 19122 56306
rect 19742 56254 19794 56306
rect 21422 56254 21474 56306
rect 22430 56254 22482 56306
rect 27134 56254 27186 56306
rect 28366 56254 28418 56306
rect 29822 56254 29874 56306
rect 31838 56254 31890 56306
rect 33182 56254 33234 56306
rect 33854 56254 33906 56306
rect 37102 56254 37154 56306
rect 37774 56254 37826 56306
rect 38558 56254 38610 56306
rect 39230 56254 39282 56306
rect 41022 56254 41074 56306
rect 41694 56254 41746 56306
rect 43934 56254 43986 56306
rect 45502 56254 45554 56306
rect 47966 56254 48018 56306
rect 48862 56254 48914 56306
rect 49534 56254 49586 56306
rect 1822 56142 1874 56194
rect 3054 56142 3106 56194
rect 5854 56142 5906 56194
rect 46062 56142 46114 56194
rect 54910 56142 54962 56194
rect 4174 56030 4226 56082
rect 12798 56030 12850 56082
rect 15038 56030 15090 56082
rect 56814 56030 56866 56082
rect 7198 55918 7250 55970
rect 12014 55918 12066 55970
rect 47182 55918 47234 55970
rect 54014 55918 54066 55970
rect 55918 55918 55970 55970
rect 57374 55918 57426 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 5742 55358 5794 55410
rect 46286 55358 46338 55410
rect 48414 55358 48466 55410
rect 55134 55358 55186 55410
rect 3054 55246 3106 55298
rect 45614 55246 45666 55298
rect 1934 55134 1986 55186
rect 3614 55134 3666 55186
rect 4286 55134 4338 55186
rect 13694 55134 13746 55186
rect 56254 55134 56306 55186
rect 57374 55134 57426 55186
rect 57934 55134 57986 55186
rect 4846 55022 4898 55074
rect 48862 55022 48914 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 2494 54686 2546 54738
rect 3166 54686 3218 54738
rect 56702 54686 56754 54738
rect 58046 54686 58098 54738
rect 1822 54574 1874 54626
rect 52222 54574 52274 54626
rect 53566 54574 53618 54626
rect 44494 54462 44546 54514
rect 51886 54462 51938 54514
rect 52894 54462 52946 54514
rect 3726 54350 3778 54402
rect 41582 54350 41634 54402
rect 43710 54350 43762 54402
rect 44942 54350 44994 54402
rect 55694 54350 55746 54402
rect 56254 54350 56306 54402
rect 55918 54238 55970 54290
rect 56814 54238 56866 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 43934 53790 43986 53842
rect 50094 53790 50146 53842
rect 3054 53678 3106 53730
rect 44158 53678 44210 53730
rect 44718 53678 44770 53730
rect 47294 53678 47346 53730
rect 1934 53566 1986 53618
rect 47966 53566 48018 53618
rect 50542 53566 50594 53618
rect 3502 53454 3554 53506
rect 46734 53454 46786 53506
rect 58046 53454 58098 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 44270 53118 44322 53170
rect 44382 53118 44434 53170
rect 45278 53118 45330 53170
rect 1822 53006 1874 53058
rect 45502 53006 45554 53058
rect 48078 53006 48130 53058
rect 58046 53006 58098 53058
rect 44158 52894 44210 52946
rect 44718 52894 44770 52946
rect 45614 52894 45666 52946
rect 48190 52894 48242 52946
rect 53006 52894 53058 52946
rect 48638 52782 48690 52834
rect 49422 52782 49474 52834
rect 50094 52782 50146 52834
rect 52222 52782 52274 52834
rect 53454 52782 53506 52834
rect 48078 52670 48130 52722
rect 48414 52670 48466 52722
rect 48638 52670 48690 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 39902 52222 39954 52274
rect 43262 52222 43314 52274
rect 45614 52222 45666 52274
rect 53454 52222 53506 52274
rect 55582 52222 55634 52274
rect 42030 52110 42082 52162
rect 42814 52110 42866 52162
rect 44830 52110 44882 52162
rect 47966 52110 48018 52162
rect 48190 52110 48242 52162
rect 49086 52110 49138 52162
rect 56254 52110 56306 52162
rect 56814 52110 56866 52162
rect 44494 51998 44546 52050
rect 45950 51998 46002 52050
rect 47294 51998 47346 52050
rect 51326 51998 51378 52050
rect 51662 51998 51714 52050
rect 44046 51886 44098 51938
rect 44606 51886 44658 51938
rect 45502 51886 45554 51938
rect 45726 51886 45778 51938
rect 46398 51886 46450 51938
rect 48750 51886 48802 51938
rect 48974 51886 49026 51938
rect 49646 51886 49698 51938
rect 50094 51886 50146 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 41918 51550 41970 51602
rect 44494 51550 44546 51602
rect 45614 51550 45666 51602
rect 49422 51550 49474 51602
rect 53454 51550 53506 51602
rect 1822 51438 1874 51490
rect 44046 51438 44098 51490
rect 44718 51438 44770 51490
rect 44830 51438 44882 51490
rect 45838 51438 45890 51490
rect 46622 51438 46674 51490
rect 46734 51438 46786 51490
rect 49646 51438 49698 51490
rect 58046 51438 58098 51490
rect 41694 51326 41746 51378
rect 45950 51326 46002 51378
rect 46398 51326 46450 51378
rect 48078 51326 48130 51378
rect 49758 51326 49810 51378
rect 48190 51214 48242 51266
rect 50206 51214 50258 51266
rect 50654 51214 50706 51266
rect 51326 51214 51378 51266
rect 52558 51214 52610 51266
rect 53006 51214 53058 51266
rect 54798 51214 54850 51266
rect 47630 51102 47682 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 49198 50766 49250 50818
rect 49870 50766 49922 50818
rect 39566 50654 39618 50706
rect 42926 50654 42978 50706
rect 46286 50654 46338 50706
rect 47630 50654 47682 50706
rect 49870 50654 49922 50706
rect 51774 50654 51826 50706
rect 55134 50654 55186 50706
rect 57262 50654 57314 50706
rect 42478 50542 42530 50594
rect 46398 50542 46450 50594
rect 47854 50542 47906 50594
rect 51438 50542 51490 50594
rect 52222 50542 52274 50594
rect 57934 50542 57986 50594
rect 41694 50430 41746 50482
rect 44718 50430 44770 50482
rect 45502 50430 45554 50482
rect 47182 50430 47234 50482
rect 48974 50430 49026 50482
rect 49422 50430 49474 50482
rect 48638 50318 48690 50370
rect 48862 50318 48914 50370
rect 50318 50318 50370 50370
rect 50878 50318 50930 50370
rect 53342 50318 53394 50370
rect 53790 50318 53842 50370
rect 54350 50318 54402 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 44494 49982 44546 50034
rect 47294 49982 47346 50034
rect 47406 49982 47458 50034
rect 49422 49982 49474 50034
rect 50430 49982 50482 50034
rect 52110 49982 52162 50034
rect 53454 49982 53506 50034
rect 58046 49982 58098 50034
rect 48638 49870 48690 49922
rect 48750 49870 48802 49922
rect 52894 49870 52946 49922
rect 53006 49870 53058 49922
rect 53678 49870 53730 49922
rect 44382 49758 44434 49810
rect 44606 49758 44658 49810
rect 44942 49758 44994 49810
rect 45614 49758 45666 49810
rect 45838 49758 45890 49810
rect 47518 49758 47570 49810
rect 47630 49758 47682 49810
rect 47966 49758 48018 49810
rect 48414 49758 48466 49810
rect 50990 49758 51042 49810
rect 51550 49758 51602 49810
rect 51774 49758 51826 49810
rect 51998 49758 52050 49810
rect 52670 49758 52722 49810
rect 53790 49758 53842 49810
rect 56142 49758 56194 49810
rect 49870 49646 49922 49698
rect 51886 49646 51938 49698
rect 54238 49646 54290 49698
rect 55358 49646 55410 49698
rect 56590 49646 56642 49698
rect 45502 49534 45554 49586
rect 49310 49534 49362 49586
rect 50206 49534 50258 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 47518 49198 47570 49250
rect 48190 49198 48242 49250
rect 51102 49198 51154 49250
rect 53566 49198 53618 49250
rect 42702 49086 42754 49138
rect 48750 49086 48802 49138
rect 49198 49086 49250 49138
rect 58046 49086 58098 49138
rect 41134 48974 41186 49026
rect 43262 48974 43314 49026
rect 44158 48974 44210 49026
rect 44494 48974 44546 49026
rect 45838 48974 45890 49026
rect 46062 48974 46114 49026
rect 48526 48974 48578 49026
rect 50094 48974 50146 49026
rect 50654 48974 50706 49026
rect 51662 48974 51714 49026
rect 52558 48974 52610 49026
rect 54574 48974 54626 49026
rect 55246 48974 55298 49026
rect 41358 48862 41410 48914
rect 44718 48862 44770 48914
rect 45950 48862 46002 48914
rect 46398 48862 46450 48914
rect 46958 48862 47010 48914
rect 47406 48862 47458 48914
rect 50318 48862 50370 48914
rect 50542 48862 50594 48914
rect 52670 48862 52722 48914
rect 53678 48862 53730 48914
rect 55918 48862 55970 48914
rect 42590 48750 42642 48802
rect 42814 48750 42866 48802
rect 47518 48750 47570 48802
rect 51662 48750 51714 48802
rect 53566 48750 53618 48802
rect 54126 48750 54178 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 49870 48414 49922 48466
rect 50318 48414 50370 48466
rect 52446 48414 52498 48466
rect 52782 48414 52834 48466
rect 57374 48414 57426 48466
rect 41694 48302 41746 48354
rect 47518 48302 47570 48354
rect 48302 48302 48354 48354
rect 53566 48302 53618 48354
rect 53902 48302 53954 48354
rect 55358 48302 55410 48354
rect 58046 48302 58098 48354
rect 42366 48190 42418 48242
rect 42590 48190 42642 48242
rect 44270 48190 44322 48242
rect 44718 48190 44770 48242
rect 45838 48190 45890 48242
rect 46510 48190 46562 48242
rect 46734 48190 46786 48242
rect 47294 48190 47346 48242
rect 51774 48190 51826 48242
rect 51998 48190 52050 48242
rect 53454 48190 53506 48242
rect 54238 48190 54290 48242
rect 44830 48078 44882 48130
rect 47630 48078 47682 48130
rect 48750 48078 48802 48130
rect 49422 48078 49474 48130
rect 50990 48078 51042 48130
rect 51550 48078 51602 48130
rect 56366 48078 56418 48130
rect 48190 47966 48242 48018
rect 49422 47966 49474 48018
rect 50206 47966 50258 48018
rect 54462 47966 54514 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 42590 47630 42642 47682
rect 44270 47630 44322 47682
rect 51998 47630 52050 47682
rect 43150 47518 43202 47570
rect 45502 47518 45554 47570
rect 46398 47518 46450 47570
rect 49310 47518 49362 47570
rect 49758 47518 49810 47570
rect 50654 47518 50706 47570
rect 51102 47518 51154 47570
rect 53342 47518 53394 47570
rect 54462 47518 54514 47570
rect 55134 47518 55186 47570
rect 57262 47518 57314 47570
rect 43374 47406 43426 47458
rect 44382 47406 44434 47458
rect 46174 47406 46226 47458
rect 47406 47406 47458 47458
rect 48078 47406 48130 47458
rect 51774 47406 51826 47458
rect 53902 47406 53954 47458
rect 54126 47406 54178 47458
rect 54350 47406 54402 47458
rect 57934 47406 57986 47458
rect 47854 47294 47906 47346
rect 48862 47294 48914 47346
rect 54462 47294 54514 47346
rect 1822 47182 1874 47234
rect 44270 47182 44322 47234
rect 46958 47182 47010 47234
rect 47630 47182 47682 47234
rect 48526 47182 48578 47234
rect 48750 47182 48802 47234
rect 50206 47182 50258 47234
rect 52334 47182 52386 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 46958 46846 47010 46898
rect 48190 46846 48242 46898
rect 48302 46846 48354 46898
rect 51214 46846 51266 46898
rect 51438 46846 51490 46898
rect 51550 46846 51602 46898
rect 53678 46846 53730 46898
rect 54798 46846 54850 46898
rect 55806 46846 55858 46898
rect 56254 46846 56306 46898
rect 57486 46846 57538 46898
rect 46174 46734 46226 46786
rect 47070 46734 47122 46786
rect 52334 46734 52386 46786
rect 53006 46734 53058 46786
rect 53118 46734 53170 46786
rect 54574 46734 54626 46786
rect 58046 46734 58098 46786
rect 46510 46622 46562 46674
rect 47294 46622 47346 46674
rect 47518 46622 47570 46674
rect 48526 46622 48578 46674
rect 48750 46622 48802 46674
rect 49982 46622 50034 46674
rect 50206 46622 50258 46674
rect 50990 46622 51042 46674
rect 52222 46622 52274 46674
rect 52558 46622 52610 46674
rect 53342 46622 53394 46674
rect 55470 46622 55522 46674
rect 48414 46510 48466 46562
rect 51326 46510 51378 46562
rect 56702 46510 56754 46562
rect 49646 46398 49698 46450
rect 54910 46398 54962 46450
rect 56030 46398 56082 46450
rect 56702 46398 56754 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 50990 46062 51042 46114
rect 55022 46062 55074 46114
rect 56030 46062 56082 46114
rect 42926 45950 42978 46002
rect 47182 45950 47234 46002
rect 50094 45950 50146 46002
rect 50766 45950 50818 46002
rect 51998 45950 52050 46002
rect 54462 45950 54514 46002
rect 54910 45950 54962 46002
rect 55918 45950 55970 46002
rect 57374 45950 57426 46002
rect 47294 45838 47346 45890
rect 48190 45838 48242 45890
rect 48750 45838 48802 45890
rect 51886 45838 51938 45890
rect 52110 45838 52162 45890
rect 52334 45838 52386 45890
rect 53454 45838 53506 45890
rect 53678 45838 53730 45890
rect 42814 45726 42866 45778
rect 43150 45726 43202 45778
rect 43374 45726 43426 45778
rect 46174 45726 46226 45778
rect 48414 45726 48466 45778
rect 48638 45726 48690 45778
rect 54014 45726 54066 45778
rect 1822 45614 1874 45666
rect 2494 45614 2546 45666
rect 46286 45614 46338 45666
rect 47742 45614 47794 45666
rect 49198 45614 49250 45666
rect 49646 45614 49698 45666
rect 51326 45614 51378 45666
rect 53678 45614 53730 45666
rect 55582 45614 55634 45666
rect 58046 45614 58098 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 46286 45278 46338 45330
rect 46398 45278 46450 45330
rect 49534 45278 49586 45330
rect 50766 45278 50818 45330
rect 1822 45166 1874 45218
rect 43598 45166 43650 45218
rect 48302 45166 48354 45218
rect 55246 45166 55298 45218
rect 58046 45166 58098 45218
rect 42702 45054 42754 45106
rect 43710 45054 43762 45106
rect 44270 45054 44322 45106
rect 46510 45054 46562 45106
rect 47742 45054 47794 45106
rect 48190 45054 48242 45106
rect 51886 45054 51938 45106
rect 53454 45054 53506 45106
rect 54462 45054 54514 45106
rect 55806 45054 55858 45106
rect 56366 45054 56418 45106
rect 42030 44942 42082 44994
rect 42814 44942 42866 44994
rect 45054 44942 45106 44994
rect 46062 44942 46114 44994
rect 48526 44942 48578 44994
rect 51998 44942 52050 44994
rect 52334 44942 52386 44994
rect 53342 44942 53394 44994
rect 45614 44830 45666 44882
rect 45838 44830 45890 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 43374 44494 43426 44546
rect 43710 44494 43762 44546
rect 44718 44494 44770 44546
rect 48190 44494 48242 44546
rect 45502 44382 45554 44434
rect 47070 44382 47122 44434
rect 51438 44382 51490 44434
rect 55022 44382 55074 44434
rect 44606 44270 44658 44322
rect 45614 44270 45666 44322
rect 45950 44270 46002 44322
rect 48638 44270 48690 44322
rect 49310 44270 49362 44322
rect 49646 44270 49698 44322
rect 52446 44270 52498 44322
rect 52782 44270 52834 44322
rect 53342 44270 53394 44322
rect 53902 44270 53954 44322
rect 57934 44270 57986 44322
rect 43486 44158 43538 44210
rect 44494 44158 44546 44210
rect 48414 44158 48466 44210
rect 52222 44158 52274 44210
rect 52670 44158 52722 44210
rect 53790 44158 53842 44210
rect 57262 44158 57314 44210
rect 53566 44046 53618 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 44046 43710 44098 43762
rect 52334 43710 52386 43762
rect 45502 43598 45554 43650
rect 48750 43598 48802 43650
rect 52558 43598 52610 43650
rect 53566 43598 53618 43650
rect 57598 43598 57650 43650
rect 45726 43486 45778 43538
rect 46174 43486 46226 43538
rect 47854 43486 47906 43538
rect 48526 43486 48578 43538
rect 52670 43486 52722 43538
rect 53118 43486 53170 43538
rect 50430 43374 50482 43426
rect 50878 43374 50930 43426
rect 51326 43374 51378 43426
rect 51774 43374 51826 43426
rect 58046 43374 58098 43426
rect 52894 43262 52946 43314
rect 53454 43262 53506 43314
rect 57262 43262 57314 43314
rect 58046 43262 58098 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 50206 42926 50258 42978
rect 50990 42926 51042 42978
rect 53454 42926 53506 42978
rect 43038 42814 43090 42866
rect 46286 42814 46338 42866
rect 48526 42814 48578 42866
rect 49422 42814 49474 42866
rect 50878 42814 50930 42866
rect 56366 42814 56418 42866
rect 40126 42702 40178 42754
rect 43598 42702 43650 42754
rect 48750 42702 48802 42754
rect 49310 42702 49362 42754
rect 49534 42702 49586 42754
rect 40798 42590 40850 42642
rect 48974 42590 49026 42642
rect 49198 42590 49250 42642
rect 49982 42590 50034 42642
rect 51550 42590 51602 42642
rect 52222 42590 52274 42642
rect 53678 42590 53730 42642
rect 54238 42590 54290 42642
rect 55246 42590 55298 42642
rect 39454 42478 39506 42530
rect 46174 42478 46226 42530
rect 46398 42478 46450 42530
rect 46622 42478 46674 42530
rect 48078 42478 48130 42530
rect 48190 42478 48242 42530
rect 48302 42478 48354 42530
rect 49758 42478 49810 42530
rect 50430 42478 50482 42530
rect 51662 42478 51714 42530
rect 52334 42478 52386 42530
rect 53566 42478 53618 42530
rect 56814 42478 56866 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 52782 42142 52834 42194
rect 47742 42030 47794 42082
rect 49646 42030 49698 42082
rect 49870 42030 49922 42082
rect 51214 42030 51266 42082
rect 54238 42030 54290 42082
rect 46398 41918 46450 41970
rect 46734 41918 46786 41970
rect 48414 41918 48466 41970
rect 52446 41918 52498 41970
rect 53678 41918 53730 41970
rect 54350 41918 54402 41970
rect 46846 41806 46898 41858
rect 48638 41806 48690 41858
rect 49534 41806 49586 41858
rect 50318 41806 50370 41858
rect 50990 41806 51042 41858
rect 53902 41806 53954 41858
rect 54126 41806 54178 41858
rect 54574 41694 54626 41746
rect 54798 41694 54850 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 47406 41358 47458 41410
rect 49086 41358 49138 41410
rect 49646 41358 49698 41410
rect 50990 41358 51042 41410
rect 52334 41358 52386 41410
rect 52670 41358 52722 41410
rect 45726 41246 45778 41298
rect 50206 41246 50258 41298
rect 51550 41246 51602 41298
rect 52110 41246 52162 41298
rect 53454 41246 53506 41298
rect 53902 41246 53954 41298
rect 54686 41246 54738 41298
rect 55134 41246 55186 41298
rect 57262 41246 57314 41298
rect 46398 41134 46450 41186
rect 46622 41134 46674 41186
rect 47294 41134 47346 41186
rect 48078 41134 48130 41186
rect 48302 41134 48354 41186
rect 48414 41134 48466 41186
rect 48862 41134 48914 41186
rect 49758 41134 49810 41186
rect 51102 41134 51154 41186
rect 57934 41134 57986 41186
rect 47406 41022 47458 41074
rect 49646 41022 49698 41074
rect 50990 41022 51042 41074
rect 1822 40910 1874 40962
rect 2494 40910 2546 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 44942 40574 44994 40626
rect 46286 40574 46338 40626
rect 46734 40574 46786 40626
rect 48302 40574 48354 40626
rect 48638 40574 48690 40626
rect 50766 40574 50818 40626
rect 51326 40574 51378 40626
rect 51662 40574 51714 40626
rect 52222 40574 52274 40626
rect 1822 40462 1874 40514
rect 46958 40462 47010 40514
rect 47070 40462 47122 40514
rect 47966 40462 48018 40514
rect 48078 40462 48130 40514
rect 49646 40462 49698 40514
rect 49758 40462 49810 40514
rect 56030 40462 56082 40514
rect 58046 40462 58098 40514
rect 40910 40350 40962 40402
rect 41694 40350 41746 40402
rect 42366 40350 42418 40402
rect 49982 40350 50034 40402
rect 50318 40350 50370 40402
rect 55134 40350 55186 40402
rect 44494 40238 44546 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 47406 39678 47458 39730
rect 48414 39678 48466 39730
rect 50318 39678 50370 39730
rect 50878 39678 50930 39730
rect 49982 39566 50034 39618
rect 49422 39454 49474 39506
rect 1822 39342 1874 39394
rect 58046 39342 58098 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 49534 38894 49586 38946
rect 49758 38782 49810 38834
rect 53678 38782 53730 38834
rect 50766 38670 50818 38722
rect 52894 38670 52946 38722
rect 54238 38670 54290 38722
rect 54574 38670 54626 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 53454 38110 53506 38162
rect 56366 37998 56418 38050
rect 55582 37886 55634 37938
rect 56814 37774 56866 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 53566 37438 53618 37490
rect 54014 37326 54066 37378
rect 54350 37326 54402 37378
rect 56254 37326 56306 37378
rect 55134 37102 55186 37154
rect 57374 37102 57426 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 48302 36542 48354 36594
rect 50430 36542 50482 36594
rect 47518 36430 47570 36482
rect 50878 36430 50930 36482
rect 54910 36318 54962 36370
rect 55246 36206 55298 36258
rect 55806 36206 55858 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 1822 35758 1874 35810
rect 56142 35646 56194 35698
rect 55358 35534 55410 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 54574 34974 54626 35026
rect 55918 34974 55970 35026
rect 58046 34974 58098 35026
rect 55134 34862 55186 34914
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 1822 31502 1874 31554
rect 2494 31502 2546 31554
rect 57374 31502 57426 31554
rect 58046 31502 58098 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 58046 31054 58098 31106
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 1822 28366 1874 28418
rect 58046 28366 58098 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1822 26798 1874 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 42814 26462 42866 26514
rect 42254 26350 42306 26402
rect 42030 26238 42082 26290
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 40462 25566 40514 25618
rect 42590 25566 42642 25618
rect 43934 25566 43986 25618
rect 3054 25454 3106 25506
rect 43374 25454 43426 25506
rect 1934 25342 1986 25394
rect 3614 25230 3666 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 58046 24782 58098 24834
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 1822 23214 1874 23266
rect 56254 23214 56306 23266
rect 55134 22990 55186 23042
rect 57374 22990 57426 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 1822 22094 1874 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 1822 21646 1874 21698
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 1822 20078 1874 20130
rect 56254 20078 56306 20130
rect 54910 19854 54962 19906
rect 57374 19854 57426 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 1822 18510 1874 18562
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 1822 16942 1874 16994
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 58046 15822 58098 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 1822 15374 1874 15426
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 1822 14254 1874 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 58046 13806 58098 13858
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 1822 12686 1874 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 58046 11118 58098 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 1822 10670 1874 10722
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 1822 9550 1874 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 1822 6414 1874 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 58046 5966 58098 6018
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 1822 4846 1874 4898
rect 58046 4846 58098 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 50766 4510 50818 4562
rect 1822 4398 1874 4450
rect 12350 4398 12402 4450
rect 56254 4398 56306 4450
rect 58046 4398 58098 4450
rect 13022 4174 13074 4226
rect 55134 4174 55186 4226
rect 57374 4174 57426 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 12798 3614 12850 3666
rect 30718 3614 30770 3666
rect 50542 3502 50594 3554
rect 11566 3390 11618 3442
rect 28590 3390 28642 3442
rect 29374 3390 29426 3442
rect 49422 3390 49474 3442
rect 1822 3278 1874 3330
rect 2494 3278 2546 3330
rect 3614 3278 3666 3330
rect 4286 3278 4338 3330
rect 13582 3278 13634 3330
rect 15038 3278 15090 3330
rect 16382 3278 16434 3330
rect 19070 3278 19122 3330
rect 22430 3278 22482 3330
rect 23102 3278 23154 3330
rect 24446 3278 24498 3330
rect 33182 3278 33234 3330
rect 35198 3278 35250 3330
rect 37102 3278 37154 3330
rect 39230 3278 39282 3330
rect 39902 3278 39954 3330
rect 46622 3278 46674 3330
rect 47294 3278 47346 3330
rect 48078 3278 48130 3330
rect 51102 3278 51154 3330
rect 51774 3278 51826 3330
rect 55918 3278 55970 3330
rect 56702 3278 56754 3330
rect 57934 3278 57986 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 32398 1710 32450 1762
rect 33182 1710 33234 1762
rect 50542 1710 50594 1762
rect 51102 1710 51154 1762
rect 55918 1710 55970 1762
rect 56702 1710 56754 1762
<< metal2 >>
rect 616 59200 840 59800
rect 1288 59304 1512 59800
rect 1288 59200 1540 59304
rect 1960 59200 2184 59800
rect 2632 59304 2856 59800
rect 3304 59304 3528 59800
rect 2632 59200 2884 59304
rect 3304 59200 3556 59304
rect 3976 59200 4200 59800
rect 4648 59304 4872 59800
rect 5320 59304 5544 59800
rect 4648 59200 4900 59304
rect 5320 59220 5572 59304
rect 5628 59276 5908 59332
rect 5628 59220 5684 59276
rect 5320 59200 5684 59220
rect 1484 54740 1540 59200
rect 1820 56194 1876 56206
rect 1820 56142 1822 56194
rect 1874 56142 1876 56194
rect 1820 55300 1876 56142
rect 2828 56196 2884 59200
rect 3164 58436 3220 58446
rect 3052 56196 3108 56206
rect 2828 56194 3108 56196
rect 2828 56142 3054 56194
rect 3106 56142 3108 56194
rect 2828 56140 3108 56142
rect 3052 56130 3108 56140
rect 1820 55234 1876 55244
rect 3052 55300 3108 55310
rect 3052 55206 3108 55244
rect 1484 54674 1540 54684
rect 1932 55186 1988 55198
rect 1932 55134 1934 55186
rect 1986 55134 1988 55186
rect 1820 54626 1876 54638
rect 1820 54574 1822 54626
rect 1874 54574 1876 54626
rect 1820 53956 1876 54574
rect 1932 54628 1988 55134
rect 2492 54740 2548 54750
rect 2492 54646 2548 54684
rect 3164 54738 3220 58380
rect 3500 55188 3556 59200
rect 4060 57204 4116 57214
rect 4060 55468 4116 57148
rect 4844 56306 4900 59200
rect 5516 59164 5684 59200
rect 4844 56254 4846 56306
rect 4898 56254 4900 56306
rect 4844 56242 4900 56254
rect 5852 56194 5908 59276
rect 5992 59200 6216 59800
rect 6664 59200 6888 59800
rect 7336 59200 7560 59800
rect 8680 59200 8904 59800
rect 9352 59304 9576 59800
rect 9352 59200 9604 59304
rect 10024 59200 10248 59800
rect 10696 59200 10920 59800
rect 11004 59276 11284 59332
rect 11368 59304 11592 59800
rect 12040 59304 12264 59800
rect 9548 56308 9604 59200
rect 9660 56308 9716 56318
rect 9548 56306 9716 56308
rect 9548 56254 9662 56306
rect 9714 56254 9716 56306
rect 9548 56252 9716 56254
rect 9660 56242 9716 56252
rect 11004 56306 11060 59276
rect 11228 59220 11284 59276
rect 11340 59220 11592 59304
rect 11228 59200 11592 59220
rect 12012 59200 12264 59304
rect 12712 59304 12936 59800
rect 13384 59304 13608 59800
rect 14056 59304 14280 59800
rect 12712 59200 12964 59304
rect 13384 59200 13636 59304
rect 14056 59200 14308 59304
rect 14728 59200 14952 59800
rect 15400 59200 15624 59800
rect 16072 59304 16296 59800
rect 16072 59200 16324 59304
rect 17416 59200 17640 59800
rect 18088 59200 18312 59800
rect 18760 59304 18984 59800
rect 19432 59304 19656 59800
rect 18760 59200 19012 59304
rect 19432 59200 19684 59304
rect 20104 59200 20328 59800
rect 20776 59304 21000 59800
rect 20776 59220 21028 59304
rect 21084 59276 21364 59332
rect 21084 59220 21140 59276
rect 20776 59200 21140 59220
rect 11228 59164 11396 59200
rect 11004 56254 11006 56306
rect 11058 56254 11060 56306
rect 11004 56242 11060 56254
rect 5852 56142 5854 56194
rect 5906 56142 5908 56194
rect 4172 56084 4228 56094
rect 4172 56082 4900 56084
rect 4172 56030 4174 56082
rect 4226 56030 4900 56082
rect 4172 56028 4900 56030
rect 4172 56018 4228 56028
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4060 55412 4340 55468
rect 3724 55300 3780 55310
rect 3612 55188 3668 55198
rect 3500 55186 3668 55188
rect 3500 55134 3614 55186
rect 3666 55134 3668 55186
rect 3500 55132 3668 55134
rect 3612 55122 3668 55132
rect 3164 54686 3166 54738
rect 3218 54686 3220 54738
rect 3164 54674 3220 54686
rect 1932 54562 1988 54572
rect 1820 53890 1876 53900
rect 3724 54402 3780 55244
rect 4284 55186 4340 55412
rect 4284 55134 4286 55186
rect 4338 55134 4340 55186
rect 4284 55122 4340 55134
rect 3724 54350 3726 54402
rect 3778 54350 3780 54402
rect 3052 53732 3108 53742
rect 3052 53730 3556 53732
rect 3052 53678 3054 53730
rect 3106 53678 3556 53730
rect 3052 53676 3556 53678
rect 3052 53666 3108 53676
rect 1932 53618 1988 53630
rect 1932 53566 1934 53618
rect 1986 53566 1988 53618
rect 1932 53284 1988 53566
rect 1932 53218 1988 53228
rect 3500 53506 3556 53676
rect 3500 53454 3502 53506
rect 3554 53454 3556 53506
rect 1820 53058 1876 53070
rect 1820 53006 1822 53058
rect 1874 53006 1876 53058
rect 1820 52612 1876 53006
rect 1820 52546 1876 52556
rect 3500 52052 3556 53454
rect 3724 52836 3780 54350
rect 4844 55074 4900 56028
rect 5740 55412 5796 55422
rect 5852 55412 5908 56142
rect 5740 55410 5908 55412
rect 5740 55358 5742 55410
rect 5794 55358 5908 55410
rect 5740 55356 5908 55358
rect 7196 55970 7252 55982
rect 7196 55918 7198 55970
rect 7250 55918 7252 55970
rect 5740 55346 5796 55356
rect 4844 55022 4846 55074
rect 4898 55022 4900 55074
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 3724 52770 3780 52780
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 3500 51986 3556 51996
rect 1820 51490 1876 51502
rect 1820 51438 1822 51490
rect 1874 51438 1876 51490
rect 1820 51268 1876 51438
rect 1820 51202 1876 51212
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4844 50708 4900 55022
rect 7196 53508 7252 55918
rect 12012 55970 12068 59200
rect 12796 56084 12852 56094
rect 12796 55990 12852 56028
rect 12012 55918 12014 55970
rect 12066 55918 12068 55970
rect 12012 55906 12068 55918
rect 12908 55188 12964 59200
rect 13580 56308 13636 59200
rect 13692 56308 13748 56318
rect 13580 56306 13748 56308
rect 13580 56254 13694 56306
rect 13746 56254 13748 56306
rect 13580 56252 13748 56254
rect 14252 56308 14308 59200
rect 14364 56308 14420 56318
rect 14252 56306 14420 56308
rect 14252 56254 14366 56306
rect 14418 56254 14420 56306
rect 14252 56252 14420 56254
rect 16268 56308 16324 59200
rect 16380 56308 16436 56318
rect 16268 56306 16436 56308
rect 16268 56254 16382 56306
rect 16434 56254 16436 56306
rect 16268 56252 16436 56254
rect 18956 56308 19012 59200
rect 19068 56308 19124 56318
rect 18956 56306 19124 56308
rect 18956 56254 19070 56306
rect 19122 56254 19124 56306
rect 18956 56252 19124 56254
rect 19628 56308 19684 59200
rect 20972 59164 21140 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19740 56308 19796 56318
rect 19628 56306 19796 56308
rect 19628 56254 19742 56306
rect 19794 56254 19796 56306
rect 19628 56252 19796 56254
rect 21308 56308 21364 59276
rect 21448 59200 21672 59800
rect 22120 59304 22344 59800
rect 22120 59200 22372 59304
rect 22792 59200 23016 59800
rect 23464 59200 23688 59800
rect 24136 59200 24360 59800
rect 24808 59200 25032 59800
rect 26152 59200 26376 59800
rect 26824 59304 27048 59800
rect 26824 59200 27076 59304
rect 27496 59200 27720 59800
rect 28168 59304 28392 59800
rect 28168 59200 28420 59304
rect 28840 59200 29064 59800
rect 29512 59304 29736 59800
rect 29512 59200 29764 59304
rect 30184 59200 30408 59800
rect 30856 59200 31080 59800
rect 31528 59304 31752 59800
rect 31528 59200 31780 59304
rect 32200 59200 32424 59800
rect 32872 59304 33096 59800
rect 33544 59304 33768 59800
rect 32872 59200 33124 59304
rect 33544 59200 33796 59304
rect 34888 59200 35112 59800
rect 35560 59200 35784 59800
rect 36232 59304 36456 59800
rect 36904 59304 37128 59800
rect 36232 59200 36484 59304
rect 36904 59200 37156 59304
rect 37576 59200 37800 59800
rect 38248 59304 38472 59800
rect 38920 59304 39144 59800
rect 38248 59200 38500 59304
rect 38920 59200 39172 59304
rect 39592 59200 39816 59800
rect 40264 59304 40488 59800
rect 40936 59304 41160 59800
rect 40264 59200 40516 59304
rect 40936 59200 41188 59304
rect 41608 59200 41832 59800
rect 42280 59200 42504 59800
rect 43624 59304 43848 59800
rect 43624 59200 43876 59304
rect 44296 59200 44520 59800
rect 44968 59200 45192 59800
rect 45640 59304 45864 59800
rect 45612 59200 45864 59304
rect 46312 59304 46536 59800
rect 46312 59200 46564 59304
rect 46984 59200 47208 59800
rect 47656 59200 47880 59800
rect 48328 59304 48552 59800
rect 49000 59304 49224 59800
rect 48328 59200 48580 59304
rect 49000 59220 49252 59304
rect 49308 59276 49588 59332
rect 49308 59220 49364 59276
rect 49000 59200 49364 59220
rect 21420 56308 21476 56318
rect 21308 56306 21476 56308
rect 21308 56254 21422 56306
rect 21474 56254 21476 56306
rect 21308 56252 21476 56254
rect 22316 56308 22372 59200
rect 22428 56308 22484 56318
rect 22316 56306 22484 56308
rect 22316 56254 22430 56306
rect 22482 56254 22484 56306
rect 22316 56252 22484 56254
rect 27020 56308 27076 59200
rect 27132 56308 27188 56318
rect 27020 56306 27188 56308
rect 27020 56254 27134 56306
rect 27186 56254 27188 56306
rect 27020 56252 27188 56254
rect 13692 56242 13748 56252
rect 14364 56242 14420 56252
rect 16380 56242 16436 56252
rect 19068 56242 19124 56252
rect 19740 56242 19796 56252
rect 21420 56242 21476 56252
rect 22428 56242 22484 56252
rect 27132 56242 27188 56252
rect 28364 56306 28420 59200
rect 28364 56254 28366 56306
rect 28418 56254 28420 56306
rect 28364 56242 28420 56254
rect 29708 56308 29764 59200
rect 29820 56308 29876 56318
rect 29708 56306 29876 56308
rect 29708 56254 29822 56306
rect 29874 56254 29876 56306
rect 29708 56252 29876 56254
rect 31724 56308 31780 59200
rect 31836 56308 31892 56318
rect 31724 56306 31892 56308
rect 31724 56254 31838 56306
rect 31890 56254 31892 56306
rect 31724 56252 31892 56254
rect 33068 56308 33124 59200
rect 33180 56308 33236 56318
rect 33068 56306 33236 56308
rect 33068 56254 33182 56306
rect 33234 56254 33236 56306
rect 33068 56252 33236 56254
rect 33740 56308 33796 59200
rect 33852 56308 33908 56318
rect 33740 56306 33908 56308
rect 33740 56254 33854 56306
rect 33906 56254 33908 56306
rect 33740 56252 33908 56254
rect 29820 56242 29876 56252
rect 31836 56242 31892 56252
rect 33180 56242 33236 56252
rect 33852 56242 33908 56252
rect 36428 56308 36484 59200
rect 37100 56642 37156 59200
rect 37100 56590 37102 56642
rect 37154 56590 37156 56642
rect 37100 56578 37156 56590
rect 37772 56642 37828 56654
rect 37772 56590 37774 56642
rect 37826 56590 37828 56642
rect 36428 56242 36484 56252
rect 37100 56308 37156 56318
rect 37100 56214 37156 56252
rect 37772 56306 37828 56590
rect 37772 56254 37774 56306
rect 37826 56254 37828 56306
rect 37772 56242 37828 56254
rect 38444 56308 38500 59200
rect 38556 56308 38612 56318
rect 38444 56306 38612 56308
rect 38444 56254 38558 56306
rect 38610 56254 38612 56306
rect 38444 56252 38612 56254
rect 39116 56308 39172 59200
rect 40460 56754 40516 59200
rect 40460 56702 40462 56754
rect 40514 56702 40516 56754
rect 40460 56690 40516 56702
rect 41020 56754 41076 56766
rect 41020 56702 41022 56754
rect 41074 56702 41076 56754
rect 39228 56308 39284 56318
rect 39116 56306 39284 56308
rect 39116 56254 39230 56306
rect 39282 56254 39284 56306
rect 39116 56252 39284 56254
rect 38556 56242 38612 56252
rect 39228 56242 39284 56252
rect 41020 56306 41076 56702
rect 41132 56642 41188 59200
rect 41132 56590 41134 56642
rect 41186 56590 41188 56642
rect 41132 56578 41188 56590
rect 41692 56642 41748 56654
rect 41692 56590 41694 56642
rect 41746 56590 41748 56642
rect 41020 56254 41022 56306
rect 41074 56254 41076 56306
rect 41020 56242 41076 56254
rect 41692 56306 41748 56590
rect 41692 56254 41694 56306
rect 41746 56254 41748 56306
rect 41692 56242 41748 56254
rect 43820 56308 43876 59200
rect 43932 56308 43988 56318
rect 43820 56306 43988 56308
rect 43820 56254 43934 56306
rect 43986 56254 43988 56306
rect 43820 56252 43988 56254
rect 43932 56242 43988 56252
rect 45500 56308 45556 56318
rect 45612 56308 45668 59200
rect 45500 56306 45668 56308
rect 45500 56254 45502 56306
rect 45554 56254 45668 56306
rect 45500 56252 45668 56254
rect 45500 56242 45556 56252
rect 45612 56196 45668 56252
rect 46508 56308 46564 59200
rect 46508 56242 46564 56252
rect 47964 56308 48020 56318
rect 48524 56308 48580 59200
rect 49196 59164 49364 59200
rect 48860 56308 48916 56318
rect 48524 56306 48916 56308
rect 48524 56254 48862 56306
rect 48914 56254 48916 56306
rect 48524 56252 48916 56254
rect 47964 56214 48020 56252
rect 48860 56242 48916 56252
rect 49532 56306 49588 59276
rect 49672 59200 49896 59800
rect 50344 59200 50568 59800
rect 51016 59200 51240 59800
rect 52360 59200 52584 59800
rect 53032 59200 53256 59800
rect 53704 59200 53928 59800
rect 54376 59200 54600 59800
rect 55048 59200 55272 59800
rect 55720 59200 55944 59800
rect 56392 59304 56616 59800
rect 56392 59200 56644 59304
rect 57064 59200 57288 59800
rect 57736 59304 57960 59800
rect 58408 59304 58632 59800
rect 59080 59304 59304 59800
rect 59752 59304 59976 59800
rect 57736 59200 57988 59304
rect 56588 56644 56644 59200
rect 57484 58436 57540 58446
rect 56588 56578 56644 56588
rect 57372 56644 57428 56654
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49532 56254 49534 56306
rect 49586 56254 49588 56306
rect 49532 56242 49588 56254
rect 46060 56196 46116 56206
rect 45612 56194 46116 56196
rect 45612 56142 46062 56194
rect 46114 56142 46116 56194
rect 45612 56140 46116 56142
rect 46060 56130 46116 56140
rect 54908 56194 54964 56206
rect 54908 56142 54910 56194
rect 54962 56142 54964 56194
rect 15036 56084 15092 56094
rect 12908 55122 12964 55132
rect 13692 55188 13748 55198
rect 13692 55094 13748 55132
rect 15036 54404 15092 56028
rect 46284 55972 46340 55982
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 46284 55410 46340 55916
rect 47180 55972 47236 55982
rect 47180 55878 47236 55916
rect 54012 55970 54068 55982
rect 54012 55918 54014 55970
rect 54066 55918 54068 55970
rect 46284 55358 46286 55410
rect 46338 55358 46340 55410
rect 46284 55346 46340 55358
rect 48412 55412 48468 55422
rect 54012 55412 54068 55918
rect 54908 55468 54964 56142
rect 56812 56082 56868 56094
rect 56812 56030 56814 56082
rect 56866 56030 56868 56082
rect 55916 55972 55972 55982
rect 55916 55878 55972 55916
rect 54908 55412 55076 55468
rect 48412 55410 48580 55412
rect 48412 55358 48414 55410
rect 48466 55358 48580 55410
rect 48412 55356 48580 55358
rect 48412 55346 48468 55356
rect 45612 55298 45668 55310
rect 45612 55246 45614 55298
rect 45666 55246 45668 55298
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 44492 54514 44548 54526
rect 44492 54462 44494 54514
rect 44546 54462 44548 54514
rect 15036 54338 15092 54348
rect 41580 54404 41636 54414
rect 41580 54310 41636 54348
rect 43708 54404 43764 54414
rect 44492 54404 44548 54462
rect 43708 54402 44324 54404
rect 43708 54350 43710 54402
rect 43762 54350 44324 54402
rect 43708 54348 44324 54350
rect 43708 54338 43764 54348
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 7196 53442 7252 53452
rect 43932 53842 43988 53854
rect 43932 53790 43934 53842
rect 43986 53790 43988 53842
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 43932 52948 43988 53790
rect 44156 53730 44212 53742
rect 44156 53678 44158 53730
rect 44210 53678 44212 53730
rect 44156 53172 44212 53678
rect 44156 53106 44212 53116
rect 44268 53170 44324 54348
rect 44268 53118 44270 53170
rect 44322 53118 44324 53170
rect 44268 53106 44324 53118
rect 44380 53172 44436 53182
rect 44380 53078 44436 53116
rect 44156 52948 44212 52958
rect 43932 52946 44212 52948
rect 43932 52894 44158 52946
rect 44210 52894 44212 52946
rect 43932 52892 44212 52894
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 39900 52274 39956 52286
rect 39900 52222 39902 52274
rect 39954 52222 39956 52274
rect 39900 52052 39956 52222
rect 42812 52276 42868 52286
rect 42028 52164 42084 52174
rect 39900 51986 39956 51996
rect 41916 52162 42084 52164
rect 41916 52110 42030 52162
rect 42082 52110 42084 52162
rect 41916 52108 42084 52110
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 41916 51602 41972 52108
rect 42028 52098 42084 52108
rect 42812 52162 42868 52220
rect 43260 52276 43316 52286
rect 43260 52182 43316 52220
rect 42812 52110 42814 52162
rect 42866 52110 42868 52162
rect 41916 51550 41918 51602
rect 41970 51550 41972 51602
rect 41916 51538 41972 51550
rect 41692 51378 41748 51390
rect 41692 51326 41694 51378
rect 41746 51326 41748 51378
rect 41692 51044 41748 51326
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 41692 50978 41748 50988
rect 35196 50922 35460 50932
rect 4844 50642 4900 50652
rect 39564 50708 39620 50718
rect 42812 50708 42868 52110
rect 44044 51940 44100 51950
rect 44044 51846 44100 51884
rect 44044 51492 44100 51502
rect 44044 51398 44100 51436
rect 42924 50708 42980 50718
rect 39564 50614 39620 50652
rect 42476 50706 42980 50708
rect 42476 50654 42926 50706
rect 42978 50654 42980 50706
rect 42476 50652 42980 50654
rect 42476 50594 42532 50652
rect 42924 50642 42980 50652
rect 42476 50542 42478 50594
rect 42530 50542 42532 50594
rect 42476 50530 42532 50542
rect 41692 50484 41748 50494
rect 41356 50482 41748 50484
rect 41356 50430 41694 50482
rect 41746 50430 41748 50482
rect 41356 50428 41748 50430
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 41132 49028 41188 49038
rect 41132 49026 41300 49028
rect 41132 48974 41134 49026
rect 41186 48974 41300 49026
rect 41132 48972 41300 48974
rect 41132 48962 41188 48972
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 41244 48468 41300 48972
rect 41356 48914 41412 50428
rect 41692 50418 41748 50428
rect 44156 50036 44212 52892
rect 44492 52276 44548 54348
rect 44940 54404 44996 54414
rect 44940 54310 44996 54348
rect 45612 54404 45668 55246
rect 45612 53844 45668 54348
rect 45612 53778 45668 53788
rect 47292 53844 47348 53854
rect 44716 53732 44772 53742
rect 44716 53638 44772 53676
rect 47292 53730 47348 53788
rect 47292 53678 47294 53730
rect 47346 53678 47348 53730
rect 47292 53620 47348 53678
rect 47292 53554 47348 53564
rect 47964 53618 48020 53630
rect 47964 53566 47966 53618
rect 48018 53566 48020 53618
rect 46732 53508 46788 53518
rect 46732 53414 46788 53452
rect 47964 53508 48020 53566
rect 47964 53442 48020 53452
rect 45276 53172 45332 53182
rect 45276 53078 45332 53116
rect 44828 53060 44884 53070
rect 44716 52948 44772 52958
rect 44716 52854 44772 52892
rect 44492 52210 44548 52220
rect 44828 52162 44884 53004
rect 45500 53060 45556 53070
rect 45500 52966 45556 53004
rect 48076 53060 48132 53070
rect 48076 52966 48132 53004
rect 45612 52948 45668 52958
rect 45612 52274 45668 52892
rect 48188 52946 48244 52958
rect 48188 52894 48190 52946
rect 48242 52894 48244 52946
rect 45612 52222 45614 52274
rect 45666 52222 45668 52274
rect 45612 52210 45668 52222
rect 48076 52722 48132 52734
rect 48076 52670 48078 52722
rect 48130 52670 48132 52722
rect 44828 52110 44830 52162
rect 44882 52110 44884 52162
rect 44828 52098 44884 52110
rect 47964 52162 48020 52174
rect 47964 52110 47966 52162
rect 48018 52110 48020 52162
rect 44492 52050 44548 52062
rect 44492 51998 44494 52050
rect 44546 51998 44548 52050
rect 44492 51602 44548 51998
rect 45948 52050 46004 52062
rect 45948 51998 45950 52050
rect 46002 51998 46004 52050
rect 44492 51550 44494 51602
rect 44546 51550 44548 51602
rect 44492 51538 44548 51550
rect 44604 51938 44660 51950
rect 44604 51886 44606 51938
rect 44658 51886 44660 51938
rect 44604 51380 44660 51886
rect 44604 51314 44660 51324
rect 44716 51940 44772 51950
rect 45500 51940 45556 51950
rect 44716 51490 44772 51884
rect 45388 51938 45556 51940
rect 45388 51886 45502 51938
rect 45554 51886 45556 51938
rect 45388 51884 45556 51886
rect 44716 51438 44718 51490
rect 44770 51438 44772 51490
rect 44716 50484 44772 51438
rect 44828 51828 44884 51838
rect 44828 51492 44884 51772
rect 44828 51360 44884 51436
rect 45388 50596 45444 51884
rect 45500 51874 45556 51884
rect 45724 51940 45780 51950
rect 45724 51846 45780 51884
rect 45948 51716 46004 51998
rect 46732 52052 46788 52062
rect 45612 51660 46004 51716
rect 46396 51940 46452 51950
rect 46396 51716 46452 51884
rect 45612 51602 45668 51660
rect 46396 51650 46452 51660
rect 45612 51550 45614 51602
rect 45666 51550 45668 51602
rect 45612 51538 45668 51550
rect 45836 51492 45892 51502
rect 46620 51492 46676 51502
rect 45836 51398 45892 51436
rect 46508 51490 46676 51492
rect 46508 51438 46622 51490
rect 46674 51438 46676 51490
rect 46508 51436 46676 51438
rect 45948 51380 46004 51390
rect 45948 51286 46004 51324
rect 46396 51380 46452 51390
rect 46396 51286 46452 51324
rect 46284 50708 46340 50718
rect 46284 50614 46340 50652
rect 44716 50390 44772 50428
rect 45276 50484 45332 50494
rect 45388 50484 45444 50540
rect 46396 50596 46452 50606
rect 46508 50596 46564 51436
rect 46620 51426 46676 51436
rect 46732 51490 46788 51996
rect 47292 52052 47348 52062
rect 47292 51958 47348 51996
rect 46732 51438 46734 51490
rect 46786 51438 46788 51490
rect 46732 50708 46788 51438
rect 46732 50642 46788 50652
rect 47628 51154 47684 51166
rect 47628 51102 47630 51154
rect 47682 51102 47684 51154
rect 47628 50706 47684 51102
rect 47628 50654 47630 50706
rect 47682 50654 47684 50706
rect 46396 50594 46564 50596
rect 46396 50542 46398 50594
rect 46450 50542 46564 50594
rect 46396 50540 46564 50542
rect 45332 50428 45444 50484
rect 45500 50482 45556 50494
rect 45500 50430 45502 50482
rect 45554 50430 45556 50482
rect 44492 50036 44548 50046
rect 44156 50034 44548 50036
rect 44156 49982 44494 50034
rect 44546 49982 44548 50034
rect 44156 49980 44548 49982
rect 44492 49970 44548 49980
rect 44268 49812 44324 49822
rect 42700 49140 42756 49150
rect 42700 49046 42756 49084
rect 44268 49140 44324 49756
rect 44380 49810 44436 49822
rect 44380 49758 44382 49810
rect 44434 49758 44436 49810
rect 44380 49252 44436 49758
rect 44604 49812 44660 49822
rect 44604 49718 44660 49756
rect 44940 49812 44996 49822
rect 44940 49718 44996 49756
rect 44380 49196 44660 49252
rect 41356 48862 41358 48914
rect 41410 48862 41412 48914
rect 41356 48850 41412 48862
rect 43260 49026 43316 49038
rect 43260 48974 43262 49026
rect 43314 48974 43316 49026
rect 42588 48802 42644 48814
rect 42588 48750 42590 48802
rect 42642 48750 42644 48802
rect 41244 48412 41748 48468
rect 41692 48354 41748 48412
rect 41692 48302 41694 48354
rect 41746 48302 41748 48354
rect 41692 48290 41748 48302
rect 42364 48242 42420 48254
rect 42364 48190 42366 48242
rect 42418 48190 42420 48242
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 42364 47460 42420 48190
rect 42588 48242 42644 48750
rect 42588 48190 42590 48242
rect 42642 48190 42644 48242
rect 42588 47682 42644 48190
rect 42588 47630 42590 47682
rect 42642 47630 42644 47682
rect 42588 47618 42644 47630
rect 42812 48802 42868 48814
rect 42812 48750 42814 48802
rect 42866 48750 42868 48802
rect 42812 47460 42868 48750
rect 43260 47684 43316 48974
rect 44156 49026 44212 49038
rect 44156 48974 44158 49026
rect 44210 48974 44212 49026
rect 44156 48916 44212 48974
rect 44156 48850 44212 48860
rect 44268 48242 44324 49084
rect 44492 49028 44548 49038
rect 44492 48934 44548 48972
rect 44604 48916 44660 49196
rect 44716 48916 44772 48926
rect 44604 48914 44772 48916
rect 44604 48862 44718 48914
rect 44770 48862 44772 48914
rect 44604 48860 44772 48862
rect 44268 48190 44270 48242
rect 44322 48190 44324 48242
rect 44268 48178 44324 48190
rect 44716 48242 44772 48860
rect 44716 48190 44718 48242
rect 44770 48190 44772 48242
rect 44716 48178 44772 48190
rect 44828 48130 44884 48142
rect 44828 48078 44830 48130
rect 44882 48078 44884 48130
rect 43260 47618 43316 47628
rect 44268 47684 44324 47694
rect 44268 47590 44324 47628
rect 43148 47572 43204 47582
rect 43148 47478 43204 47516
rect 44380 47572 44436 47582
rect 42364 47404 42868 47460
rect 43372 47458 43428 47470
rect 43372 47406 43374 47458
rect 43426 47406 43428 47458
rect 1820 47236 1876 47246
rect 1820 47142 1876 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 42364 46004 42420 47404
rect 43372 47236 43428 47406
rect 44380 47458 44436 47516
rect 44380 47406 44382 47458
rect 44434 47406 44436 47458
rect 44380 47394 44436 47406
rect 43372 47170 43428 47180
rect 44268 47236 44324 47246
rect 44268 47142 44324 47180
rect 43036 46676 43092 46686
rect 42924 46004 42980 46014
rect 42364 46002 42980 46004
rect 42364 45950 42926 46002
rect 42978 45950 42980 46002
rect 42364 45948 42980 45950
rect 42924 45938 42980 45948
rect 42700 45780 42756 45790
rect 1820 45668 1876 45678
rect 1708 45666 1876 45668
rect 1708 45614 1822 45666
rect 1874 45614 1876 45666
rect 1708 45612 1876 45614
rect 1708 45220 1764 45612
rect 1820 45602 1876 45612
rect 2492 45668 2548 45678
rect 2492 45574 2548 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 1708 45154 1764 45164
rect 1820 45218 1876 45230
rect 1820 45166 1822 45218
rect 1874 45166 1876 45218
rect 1820 44548 1876 45166
rect 42700 45106 42756 45724
rect 42700 45054 42702 45106
rect 42754 45054 42756 45106
rect 42700 45042 42756 45054
rect 42812 45778 42868 45790
rect 42812 45726 42814 45778
rect 42866 45726 42868 45778
rect 42812 45220 42868 45726
rect 42028 44994 42084 45006
rect 42028 44942 42030 44994
rect 42082 44942 42084 44994
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 1820 44482 1876 44492
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 42028 43708 42084 44942
rect 42812 44994 42868 45164
rect 42812 44942 42814 44994
rect 42866 44942 42868 44994
rect 42812 44930 42868 44942
rect 42028 43652 42868 43708
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 40124 42756 40180 42766
rect 40124 42662 40180 42700
rect 42028 42756 42084 42766
rect 39452 42644 39508 42654
rect 39452 42530 39508 42588
rect 40796 42644 40852 42654
rect 40796 42550 40852 42588
rect 39452 42478 39454 42530
rect 39506 42478 39508 42530
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 1820 40964 1876 40974
rect 1708 40962 1876 40964
rect 1708 40910 1822 40962
rect 1874 40910 1876 40962
rect 1708 40908 1876 40910
rect 1708 40516 1764 40908
rect 1820 40898 1876 40908
rect 2492 40964 2548 40974
rect 2492 40870 2548 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 1708 40450 1764 40460
rect 1820 40514 1876 40526
rect 1820 40462 1822 40514
rect 1874 40462 1876 40514
rect 1820 39844 1876 40462
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 1820 39778 1876 39788
rect 1820 39394 1876 39406
rect 1820 39342 1822 39394
rect 1874 39342 1876 39394
rect 1820 39172 1876 39342
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 1820 39106 1876 39116
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 1820 35810 1876 35822
rect 1820 35758 1822 35810
rect 1874 35758 1876 35810
rect 1820 35140 1876 35758
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 1820 35074 1876 35084
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 1820 31556 1876 31566
rect 1820 31462 1876 31500
rect 2492 31554 2548 31566
rect 2492 31502 2494 31554
rect 2546 31502 2548 31554
rect 2492 31108 2548 31502
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 2492 31042 2548 31052
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 1820 28420 1876 28430
rect 1820 28326 1876 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 1820 26964 1876 26974
rect 1820 26850 1876 26908
rect 1820 26798 1822 26850
rect 1874 26798 1876 26850
rect 1820 26786 1876 26798
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 3052 25506 3108 25518
rect 3052 25454 3054 25506
rect 3106 25454 3108 25506
rect 1932 25394 1988 25406
rect 1932 25342 1934 25394
rect 1986 25342 1988 25394
rect 1932 25060 1988 25342
rect 3052 25284 3108 25454
rect 3052 25218 3108 25228
rect 3612 25284 3668 25294
rect 3612 25190 3668 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 1932 24994 1988 25004
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 1820 23266 1876 23278
rect 1820 23214 1822 23266
rect 1874 23214 1876 23266
rect 1820 23044 1876 23214
rect 1820 22978 1876 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 1820 22148 1876 22158
rect 1708 22146 1876 22148
rect 1708 22094 1822 22146
rect 1874 22094 1876 22146
rect 1708 22092 1876 22094
rect 1708 21700 1764 22092
rect 1820 22082 1876 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 1708 21634 1764 21644
rect 1820 21698 1876 21710
rect 1820 21646 1822 21698
rect 1874 21646 1876 21698
rect 1820 21028 1876 21646
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 1820 20962 1876 20972
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 1820 20130 1876 20142
rect 1820 20078 1822 20130
rect 1874 20078 1876 20130
rect 1820 19684 1876 20078
rect 1820 19618 1876 19628
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 1820 18562 1876 18574
rect 1820 18510 1822 18562
rect 1874 18510 1876 18562
rect 1820 18340 1876 18510
rect 1820 18274 1876 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 1820 16994 1876 17006
rect 1820 16942 1822 16994
rect 1874 16942 1876 16994
rect 1820 16324 1876 16942
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 1820 16258 1876 16268
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 1820 15426 1876 15438
rect 1820 15374 1822 15426
rect 1874 15374 1876 15426
rect 1820 14980 1876 15374
rect 1820 14914 1876 14924
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 1820 14308 1876 14318
rect 1820 14214 1876 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 1820 12740 1876 12750
rect 1820 12646 1876 12684
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 1820 10722 1876 10734
rect 1820 10670 1822 10722
rect 1874 10670 1876 10722
rect 1820 10276 1876 10670
rect 1820 10210 1876 10220
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 1820 9604 1876 9614
rect 1820 9510 1876 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 1820 6466 1876 6478
rect 1820 6414 1822 6466
rect 1874 6414 1876 6466
rect 1820 6244 1876 6414
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 1820 6178 1876 6188
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 1820 4900 1876 4910
rect 1820 4806 1876 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 1820 4452 1876 4462
rect 12348 4452 12404 4462
rect 1820 4450 1988 4452
rect 1820 4398 1822 4450
rect 1874 4398 1988 4450
rect 1820 4396 1988 4398
rect 1820 4386 1876 4396
rect 1820 3332 1876 3342
rect 1484 3330 1876 3332
rect 1484 3278 1822 3330
rect 1874 3278 1876 3330
rect 1484 3276 1876 3278
rect 140 1652 196 1662
rect 140 800 196 1596
rect 1484 800 1540 3276
rect 1820 3266 1876 3276
rect 1932 2212 1988 4396
rect 12236 4450 12404 4452
rect 12236 4398 12350 4450
rect 12402 4398 12404 4450
rect 12236 4396 12404 4398
rect 11564 4228 11620 4238
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 11564 3442 11620 4172
rect 11564 3390 11566 3442
rect 11618 3390 11620 3442
rect 1932 2146 1988 2156
rect 2492 3330 2548 3342
rect 3612 3332 3668 3342
rect 4284 3332 4340 3342
rect 2492 3278 2494 3330
rect 2546 3278 2548 3330
rect 2492 1652 2548 3278
rect 2492 1586 2548 1596
rect 3500 3330 3668 3332
rect 3500 3278 3614 3330
rect 3666 3278 3668 3330
rect 3500 3276 3668 3278
rect 3500 800 3556 3276
rect 3612 3266 3668 3276
rect 4172 3330 4340 3332
rect 4172 3278 4286 3330
rect 4338 3278 4340 3330
rect 4172 3276 4340 3278
rect 4172 800 4228 3276
rect 4284 3266 4340 3276
rect 11564 800 11620 3390
rect 12236 800 12292 4396
rect 12348 4386 12404 4396
rect 13020 4228 13076 4238
rect 13020 4134 13076 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 30716 3780 30772 3790
rect 12796 3668 12852 3678
rect 12796 3574 12852 3612
rect 30716 3666 30772 3724
rect 39452 3780 39508 42478
rect 40908 40404 40964 40414
rect 40460 25618 40516 25630
rect 40460 25566 40462 25618
rect 40514 25566 40516 25618
rect 40460 25284 40516 25566
rect 40460 25218 40516 25228
rect 39452 3714 39508 3724
rect 30716 3614 30718 3666
rect 30770 3614 30772 3666
rect 30716 3602 30772 3614
rect 40908 3668 40964 40348
rect 41692 40404 41748 40414
rect 42028 40404 42084 42700
rect 41692 40402 42084 40404
rect 41692 40350 41694 40402
rect 41746 40350 42084 40402
rect 41692 40348 42084 40350
rect 42364 40404 42420 40414
rect 41692 40338 41748 40348
rect 42364 40310 42420 40348
rect 42812 26514 42868 43652
rect 43036 42866 43092 46620
rect 43148 45780 43204 45790
rect 43148 45686 43204 45724
rect 43372 45778 43428 45790
rect 43372 45726 43374 45778
rect 43426 45726 43428 45778
rect 43372 44546 43428 45726
rect 43596 45220 43652 45230
rect 43596 45126 43652 45164
rect 43372 44494 43374 44546
rect 43426 44494 43428 44546
rect 43372 44482 43428 44494
rect 43708 45106 43764 45118
rect 43708 45054 43710 45106
rect 43762 45054 43764 45106
rect 43708 44546 43764 45054
rect 44268 45108 44324 45118
rect 44268 45014 44324 45052
rect 43708 44494 43710 44546
rect 43762 44494 43764 44546
rect 43708 44436 43764 44494
rect 43708 44370 43764 44380
rect 44492 44996 44548 45006
rect 43484 44212 43540 44222
rect 43484 44118 43540 44156
rect 44492 44210 44548 44940
rect 44716 44884 44772 44894
rect 44716 44546 44772 44828
rect 44716 44494 44718 44546
rect 44770 44494 44772 44546
rect 44716 44482 44772 44494
rect 44604 44324 44660 44334
rect 44604 44230 44660 44268
rect 44492 44158 44494 44210
rect 44546 44158 44548 44210
rect 44492 44146 44548 44158
rect 44044 44100 44100 44110
rect 44044 43762 44100 44044
rect 44044 43710 44046 43762
rect 44098 43710 44100 43762
rect 44044 43698 44100 43710
rect 43036 42814 43038 42866
rect 43090 42814 43092 42866
rect 43036 42802 43092 42814
rect 43596 42756 43652 42766
rect 43596 42662 43652 42700
rect 44492 40628 44548 40638
rect 44492 40290 44548 40572
rect 44492 40238 44494 40290
rect 44546 40238 44548 40290
rect 44492 40226 44548 40238
rect 44828 37492 44884 48078
rect 45052 45108 45108 45118
rect 45052 44994 45108 45052
rect 45052 44942 45054 44994
rect 45106 44942 45108 44994
rect 45052 44100 45108 44942
rect 45052 44034 45108 44044
rect 44940 42980 44996 42990
rect 44940 40626 44996 42924
rect 44940 40574 44942 40626
rect 44994 40574 44996 40626
rect 44940 40562 44996 40574
rect 45276 40628 45332 50428
rect 45500 49586 45556 50430
rect 46396 50036 46452 50540
rect 46396 49970 46452 49980
rect 47180 50482 47236 50494
rect 47180 50430 47182 50482
rect 47234 50430 47236 50482
rect 45612 49812 45668 49822
rect 45612 49718 45668 49756
rect 45836 49812 45892 49822
rect 45836 49810 46004 49812
rect 45836 49758 45838 49810
rect 45890 49758 46004 49810
rect 45836 49756 46004 49758
rect 45836 49746 45892 49756
rect 45500 49534 45502 49586
rect 45554 49534 45556 49586
rect 45500 49028 45556 49534
rect 45500 48962 45556 48972
rect 45836 49028 45892 49038
rect 45836 48934 45892 48972
rect 45948 48916 46004 49756
rect 45948 48822 46004 48860
rect 46060 49026 46116 49038
rect 46060 48974 46062 49026
rect 46114 48974 46116 49026
rect 45836 48244 45892 48254
rect 46060 48244 46116 48974
rect 46508 49028 46564 49038
rect 46396 48914 46452 48926
rect 46396 48862 46398 48914
rect 46450 48862 46452 48914
rect 46396 48580 46452 48862
rect 46396 48514 46452 48524
rect 45836 48242 46116 48244
rect 45836 48190 45838 48242
rect 45890 48190 46116 48242
rect 45836 48188 46116 48190
rect 46396 48244 46452 48254
rect 45500 47572 45556 47582
rect 45500 47478 45556 47516
rect 45836 46900 45892 48188
rect 46396 47570 46452 48188
rect 46508 48242 46564 48972
rect 47180 49028 47236 50430
rect 47292 50484 47348 50494
rect 47292 50034 47348 50428
rect 47292 49982 47294 50034
rect 47346 49982 47348 50034
rect 47292 49970 47348 49982
rect 47404 50036 47460 50046
rect 47404 49942 47460 49980
rect 47516 49810 47572 49822
rect 47516 49758 47518 49810
rect 47570 49758 47572 49810
rect 47516 49252 47572 49758
rect 47628 49810 47684 50654
rect 47628 49758 47630 49810
rect 47682 49758 47684 49810
rect 47628 49746 47684 49758
rect 47852 50594 47908 50606
rect 47852 50542 47854 50594
rect 47906 50542 47908 50594
rect 47852 49812 47908 50542
rect 47964 50484 48020 52110
rect 48076 51378 48132 52670
rect 48188 52724 48244 52894
rect 48412 52724 48468 52734
rect 48188 52722 48468 52724
rect 48188 52670 48414 52722
rect 48466 52670 48468 52722
rect 48188 52668 48468 52670
rect 48412 52658 48468 52668
rect 48188 52164 48244 52174
rect 48188 52162 48356 52164
rect 48188 52110 48190 52162
rect 48242 52110 48356 52162
rect 48188 52108 48356 52110
rect 48188 52098 48244 52108
rect 48076 51326 48078 51378
rect 48130 51326 48132 51378
rect 48076 51314 48132 51326
rect 48188 51940 48244 51950
rect 48188 51492 48244 51884
rect 48300 51604 48356 52108
rect 48300 51538 48356 51548
rect 48188 51266 48244 51436
rect 48188 51214 48190 51266
rect 48242 51214 48244 51266
rect 48188 51202 48244 51214
rect 47964 50418 48020 50428
rect 48188 51044 48244 51054
rect 47964 49812 48020 49822
rect 47852 49756 47964 49812
rect 47964 49680 48020 49756
rect 47180 48962 47236 48972
rect 47292 49250 47572 49252
rect 47292 49198 47518 49250
rect 47570 49198 47572 49250
rect 47292 49196 47572 49198
rect 46956 48916 47012 48926
rect 46956 48822 47012 48860
rect 47180 48804 47236 48814
rect 47068 48356 47124 48366
rect 46508 48190 46510 48242
rect 46562 48190 46564 48242
rect 46508 48178 46564 48190
rect 46732 48244 46788 48254
rect 46732 48150 46788 48188
rect 46396 47518 46398 47570
rect 46450 47518 46452 47570
rect 46396 47506 46452 47518
rect 46172 47460 46228 47470
rect 46172 47366 46228 47404
rect 47068 47460 47124 48300
rect 45388 46844 45892 46900
rect 46396 47236 46452 47246
rect 46956 47236 47012 47246
rect 45388 42868 45444 46844
rect 46172 46788 46228 46798
rect 46172 46694 46228 46732
rect 46172 45778 46228 45790
rect 46172 45726 46174 45778
rect 46226 45726 46228 45778
rect 46060 44996 46116 45006
rect 46060 44902 46116 44940
rect 45612 44882 45668 44894
rect 45612 44830 45614 44882
rect 45666 44830 45668 44882
rect 45500 44436 45556 44446
rect 45500 44342 45556 44380
rect 45612 44322 45668 44830
rect 45836 44884 45892 44894
rect 45836 44790 45892 44828
rect 46172 44548 46228 45726
rect 46284 45666 46340 45678
rect 46284 45614 46286 45666
rect 46338 45614 46340 45666
rect 46284 45330 46340 45614
rect 46284 45278 46286 45330
rect 46338 45278 46340 45330
rect 46284 45266 46340 45278
rect 46396 45330 46452 47180
rect 46844 47234 47012 47236
rect 46844 47182 46958 47234
rect 47010 47182 47012 47234
rect 46844 47180 47012 47182
rect 46732 46788 46788 46798
rect 46508 46676 46564 46686
rect 46508 46582 46564 46620
rect 46732 45444 46788 46732
rect 46844 46676 46900 47180
rect 46956 47170 47012 47180
rect 47068 47012 47124 47404
rect 46956 46956 47124 47012
rect 46956 46898 47012 46956
rect 46956 46846 46958 46898
rect 47010 46846 47012 46898
rect 46956 46834 47012 46846
rect 47068 46788 47124 46798
rect 47180 46788 47236 48748
rect 47292 48692 47348 49196
rect 47516 49186 47572 49196
rect 48188 49250 48244 50988
rect 48524 50372 48580 55356
rect 54012 55346 54068 55356
rect 55020 55346 55076 55356
rect 55132 55410 55188 55422
rect 55132 55358 55134 55410
rect 55186 55358 55188 55410
rect 48860 55074 48916 55086
rect 48860 55022 48862 55074
rect 48914 55022 48916 55074
rect 48860 54740 48916 55022
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 48860 54674 48916 54684
rect 50540 54740 50596 54750
rect 50092 53842 50148 53854
rect 50092 53790 50094 53842
rect 50146 53790 50148 53842
rect 49420 53060 49476 53070
rect 50092 53060 50148 53790
rect 50540 53620 50596 54684
rect 52220 54628 52276 54638
rect 52220 54534 52276 54572
rect 53564 54628 53620 54638
rect 53564 54534 53620 54572
rect 51884 54514 51940 54526
rect 51884 54462 51886 54514
rect 51938 54462 51940 54514
rect 51884 53732 51940 54462
rect 52892 54516 52948 54526
rect 52892 54514 53060 54516
rect 52892 54462 52894 54514
rect 52946 54462 53060 54514
rect 52892 54460 53060 54462
rect 52892 54450 52948 54460
rect 51884 53666 51940 53676
rect 50540 53526 50596 53564
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50092 53004 50372 53060
rect 48636 52834 48692 52846
rect 48636 52782 48638 52834
rect 48690 52782 48692 52834
rect 48636 52722 48692 52782
rect 49420 52836 49476 53004
rect 50092 52836 50148 52846
rect 49420 52834 49588 52836
rect 49420 52782 49422 52834
rect 49474 52782 49588 52834
rect 49420 52780 49588 52782
rect 49420 52770 49476 52780
rect 48636 52670 48638 52722
rect 48690 52670 48692 52722
rect 48636 51716 48692 52670
rect 49084 52164 49140 52174
rect 48860 52162 49140 52164
rect 48860 52110 49086 52162
rect 49138 52110 49140 52162
rect 48860 52108 49140 52110
rect 48748 51940 48804 51950
rect 48748 51846 48804 51884
rect 48636 51650 48692 51660
rect 48748 50596 48804 50606
rect 48524 50306 48580 50316
rect 48636 50484 48692 50494
rect 48636 50370 48692 50428
rect 48636 50318 48638 50370
rect 48690 50318 48692 50370
rect 48636 50306 48692 50318
rect 48636 49922 48692 49934
rect 48636 49870 48638 49922
rect 48690 49870 48692 49922
rect 48412 49812 48468 49822
rect 48412 49718 48468 49756
rect 48636 49812 48692 49870
rect 48748 49922 48804 50540
rect 48748 49870 48750 49922
rect 48802 49870 48804 49922
rect 48748 49858 48804 49870
rect 48860 50370 48916 52108
rect 49084 52098 49140 52108
rect 48972 51940 49028 51950
rect 48972 51846 49028 51884
rect 48860 50318 48862 50370
rect 48914 50318 48916 50370
rect 48636 49746 48692 49756
rect 48860 49700 48916 50318
rect 48860 49634 48916 49644
rect 48972 51716 49028 51726
rect 48972 50484 49028 51660
rect 49420 51604 49476 51614
rect 49420 51510 49476 51548
rect 49532 51268 49588 52780
rect 50092 52742 50148 52780
rect 49644 51940 49700 51950
rect 49644 51492 49700 51884
rect 49644 51398 49700 51436
rect 50092 51938 50148 51950
rect 50092 51886 50094 51938
rect 50146 51886 50148 51938
rect 49756 51378 49812 51390
rect 49756 51326 49758 51378
rect 49810 51326 49812 51378
rect 49756 51268 49812 51326
rect 49532 51212 49700 51268
rect 49196 50818 49252 50830
rect 49196 50766 49198 50818
rect 49250 50766 49252 50818
rect 49196 50484 49252 50766
rect 48972 50482 49252 50484
rect 48972 50430 48974 50482
rect 49026 50430 49252 50482
rect 48972 50428 49252 50430
rect 49308 50596 49364 50606
rect 48188 49198 48190 49250
rect 48242 49198 48244 49250
rect 48188 49186 48244 49198
rect 48748 49140 48804 49150
rect 48748 49046 48804 49084
rect 48524 49028 48580 49038
rect 48524 48934 48580 48972
rect 47404 48916 47460 48926
rect 47404 48822 47460 48860
rect 47516 48804 47572 48814
rect 47516 48710 47572 48748
rect 47292 48636 47460 48692
rect 47292 48244 47348 48254
rect 47292 48150 47348 48188
rect 47404 47458 47460 48636
rect 47628 48580 47684 48590
rect 47516 48356 47572 48366
rect 47516 48262 47572 48300
rect 47628 48130 47684 48524
rect 48300 48356 48356 48366
rect 48300 48262 48356 48300
rect 47628 48078 47630 48130
rect 47682 48078 47684 48130
rect 47628 48066 47684 48078
rect 48748 48132 48804 48142
rect 48972 48132 49028 50428
rect 49308 50036 49364 50540
rect 49420 50484 49476 50494
rect 49420 50482 49588 50484
rect 49420 50430 49422 50482
rect 49474 50430 49588 50482
rect 49420 50428 49588 50430
rect 49420 50418 49476 50428
rect 49420 50036 49476 50046
rect 49308 50034 49476 50036
rect 49308 49982 49422 50034
rect 49474 49982 49476 50034
rect 49308 49980 49476 49982
rect 49420 49970 49476 49980
rect 49532 49812 49588 50428
rect 49532 49746 49588 49756
rect 49644 49924 49700 51212
rect 49756 50596 49812 51212
rect 49868 50818 49924 50830
rect 49868 50766 49870 50818
rect 49922 50766 49924 50818
rect 49868 50706 49924 50766
rect 49868 50654 49870 50706
rect 49922 50654 49924 50706
rect 49868 50642 49924 50654
rect 49756 50530 49812 50540
rect 50092 50372 50148 51886
rect 50204 51268 50260 51278
rect 50204 51174 50260 51212
rect 50316 50932 50372 53004
rect 53004 52946 53060 54460
rect 53004 52894 53006 52946
rect 53058 52894 53060 52946
rect 51660 52836 51716 52846
rect 51324 52052 51380 52062
rect 51324 52050 51492 52052
rect 51324 51998 51326 52050
rect 51378 51998 51492 52050
rect 51324 51996 51492 51998
rect 51324 51986 51380 51996
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50652 51492 50708 51502
rect 50652 51266 50708 51436
rect 50652 51214 50654 51266
rect 50706 51214 50708 51266
rect 50316 50876 50484 50932
rect 50316 50372 50372 50382
rect 50092 50370 50372 50372
rect 50092 50318 50318 50370
rect 50370 50318 50372 50370
rect 50092 50316 50372 50318
rect 48748 48130 49028 48132
rect 48748 48078 48750 48130
rect 48802 48078 49028 48130
rect 48748 48076 49028 48078
rect 49084 49588 49140 49598
rect 49308 49588 49364 49598
rect 49140 49586 49364 49588
rect 49140 49534 49310 49586
rect 49362 49534 49364 49586
rect 49140 49532 49364 49534
rect 48748 48066 48804 48076
rect 48188 48018 48244 48030
rect 48188 47966 48190 48018
rect 48242 47966 48244 48018
rect 47404 47406 47406 47458
rect 47458 47406 47460 47458
rect 47404 47394 47460 47406
rect 48076 47460 48132 47470
rect 48188 47460 48244 47966
rect 48076 47458 48244 47460
rect 48076 47406 48078 47458
rect 48130 47406 48244 47458
rect 48076 47404 48244 47406
rect 48076 47394 48132 47404
rect 47852 47346 47908 47358
rect 47852 47294 47854 47346
rect 47906 47294 47908 47346
rect 47124 46732 47236 46788
rect 47628 47234 47684 47246
rect 47628 47182 47630 47234
rect 47682 47182 47684 47234
rect 46956 46676 47012 46686
rect 46844 46620 46956 46676
rect 47068 46656 47124 46732
rect 47292 46676 47348 46686
rect 46956 45556 47012 46620
rect 47292 46582 47348 46620
rect 47516 46674 47572 46686
rect 47516 46622 47518 46674
rect 47570 46622 47572 46674
rect 47516 46452 47572 46622
rect 47516 46386 47572 46396
rect 47068 46340 47124 46350
rect 47068 45780 47124 46284
rect 47628 46340 47684 47182
rect 47852 47236 47908 47294
rect 48860 47346 48916 48076
rect 48860 47294 48862 47346
rect 48914 47294 48916 47346
rect 48524 47236 48580 47246
rect 47852 47234 48580 47236
rect 47852 47182 48526 47234
rect 48578 47182 48580 47234
rect 47852 47180 48580 47182
rect 48524 47170 48580 47180
rect 48748 47234 48804 47246
rect 48748 47182 48750 47234
rect 48802 47182 48804 47234
rect 48300 47012 48356 47022
rect 48188 46900 48244 46910
rect 48188 46806 48244 46844
rect 48300 46898 48356 46956
rect 48748 47012 48804 47182
rect 48748 46946 48804 46956
rect 48300 46846 48302 46898
rect 48354 46846 48356 46898
rect 48300 46834 48356 46846
rect 48524 46676 48580 46686
rect 47628 46274 47684 46284
rect 48412 46562 48468 46574
rect 48412 46510 48414 46562
rect 48466 46510 48468 46562
rect 48412 46116 48468 46510
rect 47180 46060 48468 46116
rect 47180 46002 47236 46060
rect 47180 45950 47182 46002
rect 47234 45950 47236 46002
rect 47180 45938 47236 45950
rect 47292 45892 47348 45902
rect 48188 45892 48244 45902
rect 47292 45890 47908 45892
rect 47292 45838 47294 45890
rect 47346 45838 47908 45890
rect 47292 45836 47908 45838
rect 47292 45826 47348 45836
rect 47068 45714 47124 45724
rect 47740 45666 47796 45678
rect 47740 45614 47742 45666
rect 47794 45614 47796 45666
rect 46956 45500 47124 45556
rect 46732 45378 46788 45388
rect 46396 45278 46398 45330
rect 46450 45278 46452 45330
rect 46396 45266 46452 45278
rect 45612 44270 45614 44322
rect 45666 44270 45668 44322
rect 45612 43708 45668 44270
rect 45836 44492 46228 44548
rect 46508 45108 46564 45118
rect 45836 43708 45892 44492
rect 45948 44324 46004 44334
rect 45948 44230 46004 44268
rect 46508 43708 46564 45052
rect 47068 44434 47124 45500
rect 47740 45106 47796 45614
rect 47852 45444 47908 45836
rect 48188 45556 48244 45836
rect 48412 45780 48468 45790
rect 48524 45780 48580 46620
rect 48748 46674 48804 46686
rect 48748 46622 48750 46674
rect 48802 46622 48804 46674
rect 48748 46004 48804 46622
rect 48860 46676 48916 47294
rect 48860 46610 48916 46620
rect 48748 45890 48804 45948
rect 48748 45838 48750 45890
rect 48802 45838 48804 45890
rect 48468 45724 48580 45780
rect 48636 45778 48692 45790
rect 48636 45726 48638 45778
rect 48690 45726 48692 45778
rect 48412 45686 48468 45724
rect 48636 45668 48692 45726
rect 48636 45602 48692 45612
rect 48188 45500 48468 45556
rect 47852 45388 48356 45444
rect 48300 45218 48356 45388
rect 48300 45166 48302 45218
rect 48354 45166 48356 45218
rect 48300 45154 48356 45166
rect 47740 45054 47742 45106
rect 47794 45054 47796 45106
rect 47740 45042 47796 45054
rect 48188 45108 48244 45118
rect 47068 44382 47070 44434
rect 47122 44382 47124 44434
rect 47068 44370 47124 44382
rect 47964 44996 48020 45006
rect 47964 43708 48020 44940
rect 48188 44546 48244 45052
rect 48188 44494 48190 44546
rect 48242 44494 48244 44546
rect 48188 44482 48244 44494
rect 48412 44210 48468 45500
rect 48748 45444 48804 45838
rect 48636 45388 48804 45444
rect 48972 45444 49028 45454
rect 48412 44158 48414 44210
rect 48466 44158 48468 44210
rect 48412 44146 48468 44158
rect 48524 44994 48580 45006
rect 48524 44942 48526 44994
rect 48578 44942 48580 44994
rect 48524 44884 48580 44942
rect 45500 43652 45668 43708
rect 45724 43652 45892 43708
rect 46172 43652 46564 43708
rect 47852 43652 48020 43708
rect 45500 43650 45556 43652
rect 45500 43598 45502 43650
rect 45554 43598 45556 43650
rect 45500 43586 45556 43598
rect 45388 42802 45444 42812
rect 45724 43538 45780 43652
rect 45724 43486 45726 43538
rect 45778 43486 45780 43538
rect 45724 41298 45780 43486
rect 46172 43538 46228 43652
rect 47852 43540 47908 43652
rect 46172 43486 46174 43538
rect 46226 43486 46228 43538
rect 46172 43474 46228 43486
rect 47740 43538 47908 43540
rect 47740 43486 47854 43538
rect 47906 43486 47908 43538
rect 47740 43484 47908 43486
rect 46284 42868 46340 42878
rect 46284 42774 46340 42812
rect 46172 42532 46228 42542
rect 46172 42438 46228 42476
rect 46396 42530 46452 42542
rect 46396 42478 46398 42530
rect 46450 42478 46452 42530
rect 46396 41972 46452 42478
rect 46396 41878 46452 41916
rect 46620 42530 46676 42542
rect 46620 42478 46622 42530
rect 46674 42478 46676 42530
rect 46620 41412 46676 42478
rect 46620 41346 46676 41356
rect 46732 42532 46788 42542
rect 46732 41970 46788 42476
rect 47740 42082 47796 43484
rect 47852 43474 47908 43484
rect 48524 43538 48580 44828
rect 48636 44322 48692 45388
rect 48636 44270 48638 44322
rect 48690 44270 48692 44322
rect 48636 44258 48692 44270
rect 48748 44212 48804 44222
rect 48748 43650 48804 44156
rect 48748 43598 48750 43650
rect 48802 43598 48804 43650
rect 48748 43586 48804 43598
rect 48524 43486 48526 43538
rect 48578 43486 48580 43538
rect 48524 43474 48580 43486
rect 48972 43428 49028 45388
rect 48524 42868 48580 42878
rect 48524 42774 48580 42812
rect 48748 42754 48804 42766
rect 48748 42702 48750 42754
rect 48802 42702 48804 42754
rect 47740 42030 47742 42082
rect 47794 42030 47796 42082
rect 47740 42018 47796 42030
rect 48076 42530 48132 42542
rect 48076 42478 48078 42530
rect 48130 42478 48132 42530
rect 46732 41918 46734 41970
rect 46786 41918 46788 41970
rect 45724 41246 45726 41298
rect 45778 41246 45780 41298
rect 45724 41234 45780 41246
rect 46396 41186 46452 41198
rect 46396 41134 46398 41186
rect 46450 41134 46452 41186
rect 46396 41076 46452 41134
rect 46620 41188 46676 41198
rect 46620 41094 46676 41132
rect 46396 41010 46452 41020
rect 45276 40562 45332 40572
rect 46284 40628 46340 40638
rect 46284 40534 46340 40572
rect 46732 40626 46788 41918
rect 48076 41972 48132 42478
rect 46844 41858 46900 41870
rect 46844 41806 46846 41858
rect 46898 41806 46900 41858
rect 46844 41188 46900 41806
rect 47964 41748 48020 41758
rect 47404 41412 47460 41422
rect 47404 41318 47460 41356
rect 46844 41122 46900 41132
rect 47292 41188 47348 41198
rect 47964 41188 48020 41692
rect 48076 41412 48132 41916
rect 48076 41346 48132 41356
rect 48188 42530 48244 42542
rect 48188 42478 48190 42530
rect 48242 42478 48244 42530
rect 48076 41188 48132 41198
rect 47292 41094 47348 41132
rect 47852 41186 48132 41188
rect 47852 41134 48078 41186
rect 48130 41134 48132 41186
rect 47852 41132 48132 41134
rect 47404 41076 47460 41086
rect 47404 40982 47460 41020
rect 46732 40574 46734 40626
rect 46786 40574 46788 40626
rect 46732 40562 46788 40574
rect 47068 40628 47124 40638
rect 46956 40516 47012 40526
rect 46956 40422 47012 40460
rect 47068 40514 47124 40572
rect 47068 40462 47070 40514
rect 47122 40462 47124 40514
rect 47068 40450 47124 40462
rect 47404 40516 47460 40526
rect 47404 39730 47460 40460
rect 47852 40516 47908 41132
rect 48076 41122 48132 41132
rect 48188 41076 48244 42478
rect 48300 42532 48356 42542
rect 48300 42438 48356 42476
rect 48748 42084 48804 42702
rect 48972 42642 49028 43372
rect 48972 42590 48974 42642
rect 49026 42590 49028 42642
rect 48972 42578 49028 42590
rect 49084 42308 49140 49532
rect 49308 49522 49364 49532
rect 49644 49252 49700 49868
rect 49868 49700 49924 49710
rect 49980 49700 50036 49710
rect 49868 49698 49980 49700
rect 49868 49646 49870 49698
rect 49922 49646 49980 49698
rect 49868 49644 49980 49646
rect 49868 49634 49924 49644
rect 49196 49196 49700 49252
rect 49196 49138 49252 49196
rect 49196 49086 49198 49138
rect 49250 49086 49252 49138
rect 49196 48804 49252 49086
rect 49980 49140 50036 49644
rect 50204 49586 50260 50316
rect 50316 50306 50372 50316
rect 50428 50036 50484 50876
rect 50652 50484 50708 51214
rect 50652 50418 50708 50428
rect 51324 51266 51380 51278
rect 51324 51214 51326 51266
rect 51378 51214 51380 51266
rect 50876 50372 50932 50382
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50428 50034 50708 50036
rect 50428 49982 50430 50034
rect 50482 49982 50708 50034
rect 50428 49980 50708 49982
rect 50428 49970 50484 49980
rect 50204 49534 50206 49586
rect 50258 49534 50260 49586
rect 50204 49522 50260 49534
rect 50316 49364 50372 49374
rect 50092 49140 50148 49150
rect 49980 49084 50092 49140
rect 49868 49028 49924 49038
rect 49196 48738 49252 48748
rect 49756 48916 49812 48926
rect 49420 48130 49476 48142
rect 49420 48078 49422 48130
rect 49474 48078 49476 48130
rect 49420 48020 49476 48078
rect 49308 48018 49476 48020
rect 49308 47966 49422 48018
rect 49474 47966 49476 48018
rect 49308 47964 49476 47966
rect 49308 47570 49364 47964
rect 49420 47954 49476 47964
rect 49308 47518 49310 47570
rect 49362 47518 49364 47570
rect 49308 47012 49364 47518
rect 49756 47572 49812 48860
rect 49868 48468 49924 48972
rect 49868 48336 49924 48412
rect 50092 49026 50148 49084
rect 50092 48974 50094 49026
rect 50146 48974 50148 49026
rect 49756 47478 49812 47516
rect 49980 47572 50036 47582
rect 49308 46946 49364 46956
rect 49532 47012 49588 47022
rect 49196 45780 49252 45790
rect 49196 45668 49252 45724
rect 49196 45666 49364 45668
rect 49196 45614 49198 45666
rect 49250 45614 49364 45666
rect 49196 45612 49364 45614
rect 49196 45602 49252 45612
rect 49308 44322 49364 45612
rect 49532 45330 49588 46956
rect 49980 46900 50036 47516
rect 49980 46674 50036 46844
rect 49980 46622 49982 46674
rect 50034 46622 50036 46674
rect 49980 46610 50036 46622
rect 50092 47236 50148 48974
rect 50204 48916 50260 48926
rect 50204 48468 50260 48860
rect 50316 48914 50372 49308
rect 50652 49026 50708 49980
rect 50652 48974 50654 49026
rect 50706 48974 50708 49026
rect 50652 48962 50708 48974
rect 50316 48862 50318 48914
rect 50370 48862 50372 48914
rect 50316 48692 50372 48862
rect 50540 48916 50596 48926
rect 50540 48822 50596 48860
rect 50876 48916 50932 50316
rect 50988 49812 51044 49822
rect 50988 49718 51044 49756
rect 51324 49812 51380 51214
rect 51436 50594 51492 51996
rect 51660 52050 51716 52780
rect 52220 52836 52276 52846
rect 53004 52836 53060 52894
rect 53452 52836 53508 52846
rect 53004 52834 53620 52836
rect 53004 52782 53454 52834
rect 53506 52782 53620 52834
rect 53004 52780 53620 52782
rect 52220 52742 52276 52780
rect 53452 52770 53508 52780
rect 51660 51998 51662 52050
rect 51714 51998 51716 52050
rect 51660 51986 51716 51998
rect 53452 52274 53508 52286
rect 53452 52222 53454 52274
rect 53506 52222 53508 52274
rect 53452 51602 53508 52222
rect 53564 52164 53620 52780
rect 55132 52276 55188 55358
rect 56252 55188 56308 55198
rect 56252 55094 56308 55132
rect 56700 55188 56756 55198
rect 56700 54738 56756 55132
rect 56700 54686 56702 54738
rect 56754 54686 56756 54738
rect 56700 54674 56756 54686
rect 55692 54402 55748 54414
rect 55692 54350 55694 54402
rect 55746 54350 55748 54402
rect 55692 54292 55748 54350
rect 56252 54402 56308 54414
rect 56252 54350 56254 54402
rect 56306 54350 56308 54402
rect 55916 54292 55972 54302
rect 55692 54290 55972 54292
rect 55692 54238 55918 54290
rect 55970 54238 55972 54290
rect 55692 54236 55972 54238
rect 55916 54226 55972 54236
rect 55132 52210 55188 52220
rect 55580 52276 55636 52286
rect 55580 52182 55636 52220
rect 56252 52164 56308 54350
rect 56812 54290 56868 56030
rect 56812 54238 56814 54290
rect 56866 54238 56868 54290
rect 56812 54226 56868 54238
rect 57260 55972 57316 55982
rect 56812 52164 56868 52174
rect 53564 52108 53844 52164
rect 53452 51550 53454 51602
rect 53506 51550 53508 51602
rect 52556 51266 52612 51278
rect 52556 51214 52558 51266
rect 52610 51214 52612 51266
rect 51436 50542 51438 50594
rect 51490 50542 51492 50594
rect 51436 50530 51492 50542
rect 51772 50706 51828 50718
rect 51772 50654 51774 50706
rect 51826 50654 51828 50706
rect 51772 50036 51828 50654
rect 52220 50594 52276 50606
rect 52220 50542 52222 50594
rect 52274 50542 52276 50594
rect 52108 50372 52164 50382
rect 51772 49970 51828 49980
rect 51884 50148 51940 50158
rect 51884 49924 51940 50092
rect 52108 50034 52164 50316
rect 52108 49982 52110 50034
rect 52162 49982 52164 50034
rect 52108 49970 52164 49982
rect 51884 49868 52052 49924
rect 51324 49746 51380 49756
rect 51548 49810 51604 49822
rect 51548 49758 51550 49810
rect 51602 49758 51604 49810
rect 51548 49700 51604 49758
rect 51772 49812 51828 49822
rect 51772 49718 51828 49756
rect 51996 49810 52052 49868
rect 51996 49758 51998 49810
rect 52050 49758 52052 49810
rect 51548 49634 51604 49644
rect 51884 49698 51940 49710
rect 51884 49646 51886 49698
rect 51938 49646 51940 49698
rect 51100 49252 51156 49262
rect 51100 49250 51828 49252
rect 51100 49198 51102 49250
rect 51154 49198 51828 49250
rect 51100 49196 51828 49198
rect 51100 49186 51156 49196
rect 51660 49028 51716 49066
rect 51660 48962 51716 48972
rect 50316 48636 50484 48692
rect 50316 48468 50372 48478
rect 50204 48466 50372 48468
rect 50204 48414 50318 48466
rect 50370 48414 50372 48466
rect 50204 48412 50372 48414
rect 50204 48018 50260 48412
rect 50316 48402 50372 48412
rect 50204 47966 50206 48018
rect 50258 47966 50260 48018
rect 50204 47954 50260 47966
rect 50428 48132 50484 48636
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50204 47236 50260 47246
rect 50092 47234 50260 47236
rect 50092 47182 50206 47234
rect 50258 47182 50260 47234
rect 50092 47180 50260 47182
rect 49644 46452 49700 46462
rect 49644 45892 49700 46396
rect 50092 46004 50148 47180
rect 50204 47170 50260 47180
rect 50204 47012 50260 47022
rect 50204 46674 50260 46956
rect 50204 46622 50206 46674
rect 50258 46622 50260 46674
rect 50204 46610 50260 46622
rect 50092 45910 50148 45948
rect 49644 45826 49700 45836
rect 49532 45278 49534 45330
rect 49586 45278 49588 45330
rect 49532 45266 49588 45278
rect 49644 45668 49700 45678
rect 49308 44270 49310 44322
rect 49362 44270 49364 44322
rect 49308 44258 49364 44270
rect 49644 44322 49700 45612
rect 49644 44270 49646 44322
rect 49698 44270 49700 44322
rect 49420 42868 49476 42878
rect 49420 42774 49476 42812
rect 49308 42754 49364 42766
rect 49308 42702 49310 42754
rect 49362 42702 49364 42754
rect 49196 42644 49252 42654
rect 49308 42644 49364 42702
rect 49532 42756 49588 42766
rect 49644 42756 49700 44270
rect 50428 43428 50484 48076
rect 50652 47572 50708 47582
rect 50876 47572 50932 48860
rect 51660 48804 51716 48814
rect 51436 48802 51716 48804
rect 51436 48750 51662 48802
rect 51714 48750 51716 48802
rect 51436 48748 51716 48750
rect 50988 48132 51044 48142
rect 50988 48038 51044 48076
rect 51100 47572 51156 47582
rect 50876 47570 51156 47572
rect 50876 47518 51102 47570
rect 51154 47518 51156 47570
rect 50876 47516 51156 47518
rect 50652 47478 50708 47516
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50988 47012 51044 47516
rect 51100 47506 51156 47516
rect 51212 47572 51268 47582
rect 50988 46946 51044 46956
rect 51100 46900 51156 46910
rect 50988 46676 51044 46686
rect 50876 46674 51044 46676
rect 50876 46622 50990 46674
rect 51042 46622 51044 46674
rect 50876 46620 51044 46622
rect 50764 46004 50820 46014
rect 50876 46004 50932 46620
rect 50988 46610 51044 46620
rect 50820 45948 50932 46004
rect 50764 45910 50820 45948
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50764 45332 50820 45342
rect 50876 45332 50932 45948
rect 50764 45330 50932 45332
rect 50764 45278 50766 45330
rect 50818 45278 50932 45330
rect 50764 45276 50932 45278
rect 50988 46116 51044 46126
rect 51100 46116 51156 46844
rect 51212 46898 51268 47516
rect 51436 47236 51492 48748
rect 51660 48738 51716 48748
rect 51548 48580 51604 48590
rect 51548 48130 51604 48524
rect 51548 48078 51550 48130
rect 51602 48078 51604 48130
rect 51548 47460 51604 48078
rect 51772 48242 51828 49196
rect 51772 48190 51774 48242
rect 51826 48190 51828 48242
rect 51772 48020 51828 48190
rect 51884 48244 51940 49646
rect 51996 49364 52052 49758
rect 51996 49298 52052 49308
rect 52220 49812 52276 50542
rect 52556 50148 52612 51214
rect 53004 51268 53060 51278
rect 53004 51266 53172 51268
rect 53004 51214 53006 51266
rect 53058 51214 53172 51266
rect 53004 51212 53172 51214
rect 53004 51202 53060 51212
rect 52556 50082 52612 50092
rect 53004 50260 53060 50270
rect 52892 49922 52948 49934
rect 52892 49870 52894 49922
rect 52946 49870 52948 49922
rect 52668 49812 52724 49822
rect 52220 49810 52724 49812
rect 52220 49758 52670 49810
rect 52722 49758 52724 49810
rect 52220 49756 52724 49758
rect 52220 49028 52276 49756
rect 52668 49746 52724 49756
rect 52668 49252 52724 49262
rect 52220 48962 52276 48972
rect 52556 49028 52612 49038
rect 52108 48468 52164 48478
rect 51996 48244 52052 48254
rect 51884 48242 52052 48244
rect 51884 48190 51998 48242
rect 52050 48190 52052 48242
rect 51884 48188 52052 48190
rect 51996 48178 52052 48188
rect 51772 47964 52052 48020
rect 51996 47682 52052 47964
rect 51996 47630 51998 47682
rect 52050 47630 52052 47682
rect 51996 47618 52052 47630
rect 51772 47460 51828 47470
rect 51548 47458 51828 47460
rect 51548 47406 51774 47458
rect 51826 47406 51828 47458
rect 51548 47404 51828 47406
rect 51772 47394 51828 47404
rect 51436 47180 51716 47236
rect 51212 46846 51214 46898
rect 51266 46846 51268 46898
rect 51212 46834 51268 46846
rect 51436 47012 51492 47022
rect 51436 46898 51492 46956
rect 51436 46846 51438 46898
rect 51490 46846 51492 46898
rect 51436 46834 51492 46846
rect 51548 46900 51604 46910
rect 51548 46806 51604 46844
rect 50988 46114 51156 46116
rect 50988 46062 50990 46114
rect 51042 46062 51156 46114
rect 50988 46060 51156 46062
rect 51324 46562 51380 46574
rect 51324 46510 51326 46562
rect 51378 46510 51380 46562
rect 50988 45668 51044 46060
rect 51324 45892 51380 46510
rect 51324 45826 51380 45836
rect 50764 45266 50820 45276
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50316 43426 50484 43428
rect 50316 43374 50430 43426
rect 50482 43374 50484 43426
rect 50316 43372 50484 43374
rect 50204 42978 50260 42990
rect 50204 42926 50206 42978
rect 50258 42926 50260 42978
rect 49532 42754 49700 42756
rect 49532 42702 49534 42754
rect 49586 42702 49700 42754
rect 49532 42700 49700 42702
rect 49868 42868 49924 42878
rect 49532 42690 49588 42700
rect 49196 42642 49364 42644
rect 49196 42590 49198 42642
rect 49250 42590 49364 42642
rect 49196 42588 49364 42590
rect 49196 42578 49252 42588
rect 49756 42530 49812 42542
rect 49756 42478 49758 42530
rect 49810 42478 49812 42530
rect 49756 42308 49812 42478
rect 48412 42028 48804 42084
rect 48860 42252 49812 42308
rect 48412 41970 48468 42028
rect 48412 41918 48414 41970
rect 48466 41918 48468 41970
rect 48412 41906 48468 41918
rect 48412 41300 48468 41310
rect 48300 41188 48356 41198
rect 48300 41094 48356 41132
rect 48412 41186 48468 41244
rect 48412 41134 48414 41186
rect 48466 41134 48468 41186
rect 48412 41122 48468 41134
rect 48188 41010 48244 41020
rect 47852 40450 47908 40460
rect 47964 40628 48020 40638
rect 47964 40514 48020 40572
rect 48300 40628 48356 40638
rect 48524 40628 48580 42028
rect 48636 41860 48692 41870
rect 48636 41766 48692 41804
rect 48860 41186 48916 42252
rect 49644 42084 49700 42094
rect 49084 42082 49700 42084
rect 49084 42030 49646 42082
rect 49698 42030 49700 42082
rect 49084 42028 49700 42030
rect 49084 41410 49140 42028
rect 49644 42018 49700 42028
rect 49756 41972 49812 42252
rect 49868 42082 49924 42812
rect 49868 42030 49870 42082
rect 49922 42030 49924 42082
rect 49868 42018 49924 42030
rect 49980 42642 50036 42654
rect 49980 42590 49982 42642
rect 50034 42590 50036 42642
rect 49532 41860 49588 41870
rect 49532 41766 49588 41804
rect 49084 41358 49086 41410
rect 49138 41358 49140 41410
rect 49084 41346 49140 41358
rect 49644 41412 49700 41422
rect 49644 41318 49700 41356
rect 48860 41134 48862 41186
rect 48914 41134 48916 41186
rect 48860 41122 48916 41134
rect 49756 41186 49812 41916
rect 49980 41748 50036 42590
rect 49980 41682 50036 41692
rect 49756 41134 49758 41186
rect 49810 41134 49812 41186
rect 49644 41076 49700 41086
rect 49644 40982 49700 41020
rect 49756 40740 49812 41134
rect 50204 41298 50260 42926
rect 50316 41858 50372 43372
rect 50428 43362 50484 43372
rect 50876 43428 50932 43438
rect 50876 43334 50932 43372
rect 50988 42978 51044 45612
rect 51324 45668 51380 45678
rect 51324 45574 51380 45612
rect 51436 45556 51492 45566
rect 51436 44434 51492 45500
rect 51436 44382 51438 44434
rect 51490 44382 51492 44434
rect 51436 44370 51492 44382
rect 51212 43652 51268 43662
rect 50988 42926 50990 42978
rect 51042 42926 51044 42978
rect 50876 42868 50932 42878
rect 50988 42868 51044 42926
rect 50876 42866 51044 42868
rect 50876 42814 50878 42866
rect 50930 42814 51044 42866
rect 50876 42812 51044 42814
rect 51100 43428 51156 43438
rect 50876 42802 50932 42812
rect 50428 42530 50484 42542
rect 50428 42478 50430 42530
rect 50482 42478 50484 42530
rect 50428 41972 50484 42478
rect 50988 42532 51044 42542
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50428 41906 50484 41916
rect 50316 41806 50318 41858
rect 50370 41806 50372 41858
rect 50316 41748 50372 41806
rect 50988 41858 51044 42476
rect 50988 41806 50990 41858
rect 51042 41806 51044 41858
rect 50316 41682 50372 41692
rect 50876 41748 50932 41758
rect 50204 41246 50206 41298
rect 50258 41246 50260 41298
rect 50204 41076 50260 41246
rect 50876 41076 50932 41692
rect 50988 41410 51044 41806
rect 50988 41358 50990 41410
rect 51042 41358 51044 41410
rect 50988 41346 51044 41358
rect 51100 41300 51156 43372
rect 51212 42084 51268 43596
rect 51660 43652 51716 47180
rect 51996 46676 52052 46686
rect 51884 46452 51940 46462
rect 51884 45890 51940 46396
rect 51884 45838 51886 45890
rect 51938 45838 51940 45890
rect 51884 45826 51940 45838
rect 51996 46002 52052 46620
rect 52108 46452 52164 48412
rect 52444 48468 52500 48478
rect 52556 48468 52612 48972
rect 52668 48914 52724 49196
rect 52668 48862 52670 48914
rect 52722 48862 52724 48914
rect 52668 48850 52724 48862
rect 52444 48466 52612 48468
rect 52444 48414 52446 48466
rect 52498 48414 52612 48466
rect 52444 48412 52612 48414
rect 52780 48692 52836 48702
rect 52780 48466 52836 48636
rect 52780 48414 52782 48466
rect 52834 48414 52836 48466
rect 52444 48402 52500 48412
rect 52780 47572 52836 48414
rect 52892 48468 52948 49870
rect 53004 49924 53060 50204
rect 53004 49792 53060 49868
rect 53116 49700 53172 51212
rect 53340 50372 53396 50382
rect 53340 50278 53396 50316
rect 53452 50260 53508 51550
rect 53788 51268 53844 52108
rect 56028 52162 56868 52164
rect 56028 52110 56254 52162
rect 56306 52110 56814 52162
rect 56866 52110 56868 52162
rect 56028 52108 56868 52110
rect 54796 51268 54852 51278
rect 53788 51266 54852 51268
rect 53788 51214 54798 51266
rect 54850 51214 54852 51266
rect 53788 51212 54852 51214
rect 53788 50372 53844 50382
rect 54012 50372 54068 50382
rect 54348 50372 54404 50382
rect 53788 50370 53956 50372
rect 53788 50318 53790 50370
rect 53842 50318 53956 50370
rect 53788 50316 53956 50318
rect 53788 50306 53844 50316
rect 53452 50194 53508 50204
rect 53452 50036 53508 50046
rect 53452 49942 53508 49980
rect 53676 49922 53732 49934
rect 53676 49870 53678 49922
rect 53730 49870 53732 49922
rect 53116 49634 53172 49644
rect 53452 49700 53508 49710
rect 52892 48402 52948 48412
rect 53340 48804 53396 48814
rect 52780 47506 52836 47516
rect 53340 47570 53396 48748
rect 53452 48580 53508 49644
rect 53564 49252 53620 49262
rect 53676 49252 53732 49870
rect 53620 49196 53732 49252
rect 53788 49810 53844 49822
rect 53788 49758 53790 49810
rect 53842 49758 53844 49810
rect 53564 49120 53620 49196
rect 53788 49028 53844 49758
rect 53788 48962 53844 48972
rect 53900 49812 53956 50316
rect 53676 48916 53732 48926
rect 53676 48822 53732 48860
rect 53564 48804 53620 48814
rect 53564 48710 53620 48748
rect 53900 48804 53956 49756
rect 53900 48738 53956 48748
rect 54012 49028 54068 50316
rect 53452 48242 53508 48524
rect 53788 48468 53844 48478
rect 53452 48190 53454 48242
rect 53506 48190 53508 48242
rect 53452 48178 53508 48190
rect 53564 48354 53620 48366
rect 53564 48302 53566 48354
rect 53618 48302 53620 48354
rect 53340 47518 53342 47570
rect 53394 47518 53396 47570
rect 52332 47234 52388 47246
rect 52332 47182 52334 47234
rect 52386 47182 52388 47234
rect 52332 46788 52388 47182
rect 53340 47124 53396 47518
rect 53564 48132 53620 48302
rect 53564 47348 53620 48076
rect 53788 47460 53844 48412
rect 53900 48356 53956 48366
rect 54012 48356 54068 48972
rect 54236 50370 54404 50372
rect 54236 50318 54350 50370
rect 54402 50318 54404 50370
rect 54236 50316 54404 50318
rect 54236 49698 54292 50316
rect 54348 50306 54404 50316
rect 54236 49646 54238 49698
rect 54290 49646 54292 49698
rect 53900 48354 54068 48356
rect 53900 48302 53902 48354
rect 53954 48302 54068 48354
rect 53900 48300 54068 48302
rect 53900 48290 53956 48300
rect 53900 47460 53956 47470
rect 53788 47458 53956 47460
rect 53788 47406 53902 47458
rect 53954 47406 53956 47458
rect 53788 47404 53956 47406
rect 54012 47460 54068 48300
rect 54124 48802 54180 48814
rect 54124 48750 54126 48802
rect 54178 48750 54180 48802
rect 54124 48580 54180 48750
rect 54124 47684 54180 48524
rect 54236 48468 54292 49646
rect 54572 49028 54628 49038
rect 54572 48934 54628 48972
rect 54236 48242 54292 48412
rect 54236 48190 54238 48242
rect 54290 48190 54292 48242
rect 54236 48178 54292 48190
rect 54460 48916 54516 48926
rect 54460 48018 54516 48860
rect 54796 48916 54852 51212
rect 55132 50706 55188 50718
rect 55132 50654 55134 50706
rect 55186 50654 55188 50706
rect 55132 50484 55188 50654
rect 55132 50418 55188 50428
rect 55356 49700 55412 49710
rect 55356 49606 55412 49644
rect 54796 48850 54852 48860
rect 55244 49026 55300 49038
rect 55244 48974 55246 49026
rect 55298 48974 55300 49026
rect 55244 48916 55300 48974
rect 55244 48850 55300 48860
rect 55916 48914 55972 48926
rect 55916 48862 55918 48914
rect 55970 48862 55972 48914
rect 54460 47966 54462 48018
rect 54514 47966 54516 48018
rect 54460 47908 54516 47966
rect 55356 48356 55412 48366
rect 54460 47852 54852 47908
rect 54124 47628 54404 47684
rect 54124 47460 54180 47470
rect 54012 47458 54180 47460
rect 54012 47406 54126 47458
rect 54178 47406 54180 47458
rect 54012 47404 54180 47406
rect 53900 47394 53956 47404
rect 54124 47394 54180 47404
rect 54348 47458 54404 47628
rect 54460 47572 54516 47582
rect 54460 47570 54628 47572
rect 54460 47518 54462 47570
rect 54514 47518 54628 47570
rect 54460 47516 54628 47518
rect 54460 47506 54516 47516
rect 54348 47406 54350 47458
rect 54402 47406 54404 47458
rect 53564 47282 53620 47292
rect 53340 47068 53732 47124
rect 53004 46956 53508 47012
rect 52668 46788 52724 46798
rect 52332 46786 52500 46788
rect 52332 46734 52334 46786
rect 52386 46734 52500 46786
rect 52332 46732 52500 46734
rect 52332 46722 52388 46732
rect 52220 46676 52276 46686
rect 52220 46582 52276 46620
rect 52108 46396 52276 46452
rect 51996 45950 51998 46002
rect 52050 45950 52052 46002
rect 51884 45556 51940 45566
rect 51884 45106 51940 45500
rect 51884 45054 51886 45106
rect 51938 45054 51940 45106
rect 51884 45042 51940 45054
rect 51996 44994 52052 45950
rect 52108 45890 52164 45902
rect 52108 45838 52110 45890
rect 52162 45838 52164 45890
rect 52108 45668 52164 45838
rect 52108 45602 52164 45612
rect 51996 44942 51998 44994
rect 52050 44942 52052 44994
rect 51996 44930 52052 44942
rect 52220 44436 52276 46396
rect 52332 45892 52388 45902
rect 52332 45798 52388 45836
rect 52444 45556 52500 46732
rect 52556 46676 52612 46686
rect 52668 46676 52724 46732
rect 52556 46674 52724 46676
rect 52556 46622 52558 46674
rect 52610 46622 52724 46674
rect 52556 46620 52724 46622
rect 52556 46610 52612 46620
rect 52444 45490 52500 45500
rect 52668 45892 52724 46620
rect 52332 44996 52388 45006
rect 52332 44994 52612 44996
rect 52332 44942 52334 44994
rect 52386 44942 52612 44994
rect 52332 44940 52612 44942
rect 52332 44930 52388 44940
rect 52108 44380 52276 44436
rect 52444 44548 52500 44558
rect 52108 43708 52164 44380
rect 52444 44324 52500 44492
rect 52332 44322 52500 44324
rect 52332 44270 52446 44322
rect 52498 44270 52500 44322
rect 52332 44268 52500 44270
rect 52220 44212 52276 44222
rect 52220 44118 52276 44156
rect 52220 43764 52276 43774
rect 52108 43652 52276 43708
rect 52332 43762 52388 44268
rect 52444 44258 52500 44268
rect 52556 43876 52612 44940
rect 52668 44210 52724 45836
rect 53004 46786 53060 46956
rect 53004 46734 53006 46786
rect 53058 46734 53060 46786
rect 53004 44548 53060 46734
rect 53116 46788 53172 46798
rect 53116 46694 53172 46732
rect 53340 46674 53396 46686
rect 53340 46622 53342 46674
rect 53394 46622 53396 46674
rect 53340 44994 53396 46622
rect 53452 45890 53508 46956
rect 53676 46900 53732 47068
rect 53676 46768 53732 46844
rect 54348 46004 54404 47406
rect 54460 47348 54516 47358
rect 54460 47254 54516 47292
rect 54572 46786 54628 47516
rect 54796 46898 54852 47852
rect 55132 47684 55188 47694
rect 55132 47570 55188 47628
rect 55132 47518 55134 47570
rect 55186 47518 55188 47570
rect 55132 47348 55188 47518
rect 55132 47282 55188 47292
rect 54796 46846 54798 46898
rect 54850 46846 54852 46898
rect 54796 46834 54852 46846
rect 55356 46900 55412 48300
rect 55356 46834 55412 46844
rect 55804 46900 55860 46910
rect 55916 46900 55972 48862
rect 56028 48916 56084 52108
rect 56252 52098 56308 52108
rect 56812 52098 56868 52108
rect 57260 50706 57316 55916
rect 57372 55970 57428 56588
rect 57372 55918 57374 55970
rect 57426 55918 57428 55970
rect 57372 55906 57428 55918
rect 57372 55188 57428 55198
rect 57484 55188 57540 58380
rect 57372 55186 57540 55188
rect 57372 55134 57374 55186
rect 57426 55134 57540 55186
rect 57372 55132 57540 55134
rect 57932 55186 57988 59200
rect 58380 59200 58632 59304
rect 59052 59200 59304 59304
rect 59724 59200 59976 59304
rect 57932 55134 57934 55186
rect 57986 55134 57988 55186
rect 57372 55122 57428 55132
rect 57932 55122 57988 55134
rect 58044 57428 58100 57438
rect 58044 54738 58100 57372
rect 58380 55412 58436 59200
rect 58380 55346 58436 55356
rect 59052 55188 59108 59200
rect 59724 57428 59780 59200
rect 59724 57362 59780 57372
rect 59052 55122 59108 55132
rect 58044 54686 58046 54738
rect 58098 54686 58100 54738
rect 58044 54674 58100 54686
rect 57260 50654 57262 50706
rect 57314 50654 57316 50706
rect 57260 50642 57316 50654
rect 57932 53620 57988 53630
rect 57932 50594 57988 53564
rect 58044 53506 58100 53518
rect 58044 53454 58046 53506
rect 58098 53454 58100 53506
rect 58044 53284 58100 53454
rect 58044 53218 58100 53228
rect 58044 53058 58100 53070
rect 58044 53006 58046 53058
rect 58098 53006 58100 53058
rect 58044 52612 58100 53006
rect 58044 52546 58100 52556
rect 58044 51490 58100 51502
rect 58044 51438 58046 51490
rect 58098 51438 58100 51490
rect 58044 51268 58100 51438
rect 58044 51202 58100 51212
rect 57932 50542 57934 50594
rect 57986 50542 57988 50594
rect 57932 50036 57988 50542
rect 58044 50036 58100 50046
rect 57932 50034 58100 50036
rect 57932 49982 58046 50034
rect 58098 49982 58100 50034
rect 57932 49980 58100 49982
rect 56140 49810 56196 49822
rect 56140 49758 56142 49810
rect 56194 49758 56196 49810
rect 56140 49140 56196 49758
rect 56588 49700 56644 49710
rect 56140 49074 56196 49084
rect 56252 49698 56644 49700
rect 56252 49646 56590 49698
rect 56642 49646 56644 49698
rect 56252 49644 56644 49646
rect 56140 48916 56196 48926
rect 56028 48860 56140 48916
rect 55804 46898 55972 46900
rect 55804 46846 55806 46898
rect 55858 46846 55972 46898
rect 55804 46844 55972 46846
rect 55804 46834 55860 46844
rect 54572 46734 54574 46786
rect 54626 46734 54628 46786
rect 54572 46722 54628 46734
rect 55468 46676 55524 46686
rect 55244 46674 55524 46676
rect 55244 46622 55470 46674
rect 55522 46622 55524 46674
rect 55244 46620 55524 46622
rect 54908 46452 54964 46462
rect 54908 46358 54964 46396
rect 55020 46114 55076 46126
rect 55020 46062 55022 46114
rect 55074 46062 55076 46114
rect 54460 46004 54516 46014
rect 54908 46004 54964 46014
rect 55020 46004 55076 46062
rect 54348 46002 55076 46004
rect 54348 45950 54462 46002
rect 54514 45950 54910 46002
rect 54962 45950 55076 46002
rect 54348 45948 55076 45950
rect 54460 45938 54516 45948
rect 54908 45938 54964 45948
rect 53452 45838 53454 45890
rect 53506 45838 53508 45890
rect 53452 45826 53508 45838
rect 53676 45892 53732 45930
rect 53676 45826 53732 45836
rect 54012 45778 54068 45790
rect 54012 45726 54014 45778
rect 54066 45726 54068 45778
rect 53676 45666 53732 45678
rect 53676 45614 53678 45666
rect 53730 45614 53732 45666
rect 53452 45108 53508 45118
rect 53452 45106 53620 45108
rect 53452 45054 53454 45106
rect 53506 45054 53620 45106
rect 53452 45052 53620 45054
rect 53452 45042 53508 45052
rect 53340 44942 53342 44994
rect 53394 44942 53396 44994
rect 53340 44930 53396 44942
rect 53004 44482 53060 44492
rect 52780 44324 52836 44334
rect 53340 44324 53396 44334
rect 52780 44322 53396 44324
rect 52780 44270 52782 44322
rect 52834 44270 53342 44322
rect 53394 44270 53396 44322
rect 52780 44268 53396 44270
rect 53564 44324 53620 45052
rect 53676 44436 53732 45614
rect 54012 45108 54068 45726
rect 54460 45108 54516 45118
rect 54012 45106 54516 45108
rect 54012 45054 54462 45106
rect 54514 45054 54516 45106
rect 54012 45052 54516 45054
rect 53676 44380 53956 44436
rect 53564 44268 53844 44324
rect 52780 44258 52836 44268
rect 53340 44258 53396 44268
rect 52668 44158 52670 44210
rect 52722 44158 52724 44210
rect 52668 44146 52724 44158
rect 53788 44210 53844 44268
rect 53900 44322 53956 44380
rect 53900 44270 53902 44322
rect 53954 44270 53956 44322
rect 53900 44258 53956 44270
rect 53788 44158 53790 44210
rect 53842 44158 53844 44210
rect 53564 44100 53620 44110
rect 53564 44006 53620 44044
rect 52556 43820 52724 43876
rect 52332 43710 52334 43762
rect 52386 43710 52388 43762
rect 52332 43698 52388 43710
rect 51660 43586 51716 43596
rect 51212 41952 51268 42028
rect 51324 43426 51380 43438
rect 51772 43428 51828 43438
rect 51324 43374 51326 43426
rect 51378 43374 51380 43426
rect 51324 42644 51380 43374
rect 51548 43426 51828 43428
rect 51548 43374 51774 43426
rect 51826 43374 51828 43426
rect 51548 43372 51828 43374
rect 51548 42644 51604 43372
rect 51772 43362 51828 43372
rect 51324 42642 51604 42644
rect 51324 42590 51550 42642
rect 51602 42590 51604 42642
rect 51324 42588 51604 42590
rect 51324 41972 51380 42588
rect 51548 42578 51604 42588
rect 52220 42642 52276 43652
rect 52556 43652 52612 43662
rect 52556 43558 52612 43596
rect 52668 43538 52724 43820
rect 52668 43486 52670 43538
rect 52722 43486 52724 43538
rect 52668 43428 52724 43486
rect 53116 43764 53172 43774
rect 53116 43538 53172 43708
rect 53564 43652 53620 43662
rect 53620 43596 53732 43652
rect 53564 43558 53620 43596
rect 53116 43486 53118 43538
rect 53170 43486 53172 43538
rect 53116 43474 53172 43486
rect 52220 42590 52222 42642
rect 52274 42590 52276 42642
rect 51324 41906 51380 41916
rect 51660 42530 51716 42542
rect 51660 42478 51662 42530
rect 51714 42478 51716 42530
rect 51660 41972 51716 42478
rect 51660 41906 51716 41916
rect 52108 42084 52164 42094
rect 51548 41300 51604 41310
rect 51156 41298 51604 41300
rect 51156 41246 51550 41298
rect 51602 41246 51604 41298
rect 51156 41244 51604 41246
rect 51100 41186 51156 41244
rect 51100 41134 51102 41186
rect 51154 41134 51156 41186
rect 51100 41122 51156 41134
rect 50988 41076 51044 41086
rect 50876 41074 51044 41076
rect 50876 41022 50990 41074
rect 51042 41022 51044 41074
rect 50876 41020 51044 41022
rect 50204 41010 50260 41020
rect 50988 40852 51044 41020
rect 49644 40684 49812 40740
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50988 40786 51044 40796
rect 51324 41076 51380 41086
rect 50556 40730 50820 40740
rect 48300 40626 48580 40628
rect 48300 40574 48302 40626
rect 48354 40574 48580 40626
rect 48300 40572 48580 40574
rect 48636 40628 48692 40638
rect 48300 40562 48356 40572
rect 48636 40534 48692 40572
rect 49644 40628 49700 40684
rect 47964 40462 47966 40514
rect 48018 40462 48020 40514
rect 47964 40450 48020 40462
rect 48076 40514 48132 40526
rect 48076 40462 48078 40514
rect 48130 40462 48132 40514
rect 48076 40404 48132 40462
rect 49644 40514 49700 40572
rect 50764 40628 50820 40638
rect 50820 40572 50932 40628
rect 50764 40534 50820 40572
rect 49644 40462 49646 40514
rect 49698 40462 49700 40514
rect 49644 40450 49700 40462
rect 49756 40514 49812 40526
rect 49756 40462 49758 40514
rect 49810 40462 49812 40514
rect 48076 40338 48132 40348
rect 48412 40404 48468 40414
rect 47404 39678 47406 39730
rect 47458 39678 47460 39730
rect 47404 39666 47460 39678
rect 48412 39730 48468 40348
rect 49756 40404 49812 40462
rect 49756 40338 49812 40348
rect 49980 40402 50036 40414
rect 49980 40350 49982 40402
rect 50034 40350 50036 40402
rect 48412 39678 48414 39730
rect 48466 39678 48468 39730
rect 48412 39666 48468 39678
rect 49980 39618 50036 40350
rect 50316 40404 50372 40414
rect 50316 40310 50372 40348
rect 50316 39732 50372 39742
rect 50316 39638 50372 39676
rect 50876 39730 50932 40572
rect 51324 40626 51380 41020
rect 51324 40574 51326 40626
rect 51378 40574 51380 40626
rect 51324 40562 51380 40574
rect 51548 40628 51604 41244
rect 52108 41298 52164 42028
rect 52108 41246 52110 41298
rect 52162 41246 52164 41298
rect 52108 41234 52164 41246
rect 52220 41076 52276 42590
rect 52444 43372 52948 43428
rect 52332 42530 52388 42542
rect 52332 42478 52334 42530
rect 52386 42478 52388 42530
rect 52332 41860 52388 42478
rect 52332 41794 52388 41804
rect 52444 41970 52500 43372
rect 52892 43314 52948 43372
rect 52892 43262 52894 43314
rect 52946 43262 52948 43314
rect 52892 43250 52948 43262
rect 53452 43314 53508 43326
rect 53452 43262 53454 43314
rect 53506 43262 53508 43314
rect 53452 42978 53508 43262
rect 53452 42926 53454 42978
rect 53506 42926 53508 42978
rect 53452 42914 53508 42926
rect 53452 42644 53508 42654
rect 52444 41918 52446 41970
rect 52498 41918 52500 41970
rect 52332 41412 52388 41422
rect 52444 41412 52500 41918
rect 52780 42194 52836 42206
rect 52780 42142 52782 42194
rect 52834 42142 52836 42194
rect 52780 42084 52836 42142
rect 52332 41410 52500 41412
rect 52332 41358 52334 41410
rect 52386 41358 52500 41410
rect 52332 41356 52500 41358
rect 52668 41412 52724 41422
rect 52332 41346 52388 41356
rect 52668 41318 52724 41356
rect 52220 41020 52388 41076
rect 51548 40562 51604 40572
rect 51660 40852 51716 40862
rect 51660 40626 51716 40796
rect 51660 40574 51662 40626
rect 51714 40574 51716 40626
rect 51660 40562 51716 40574
rect 52220 40628 52276 40638
rect 52220 40534 52276 40572
rect 52332 40404 52388 41020
rect 52332 40338 52388 40348
rect 50876 39678 50878 39730
rect 50930 39678 50932 39730
rect 49980 39566 49982 39618
rect 50034 39566 50036 39618
rect 49980 39554 50036 39566
rect 49420 39506 49476 39518
rect 49420 39454 49422 39506
rect 49474 39454 49476 39506
rect 49420 39172 49476 39454
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 49420 39116 49812 39172
rect 50556 39162 50820 39172
rect 44828 37426 44884 37436
rect 49532 38946 49588 38958
rect 49532 38894 49534 38946
rect 49586 38894 49588 38946
rect 48300 37268 48356 37278
rect 48300 36594 48356 37212
rect 49532 37268 49588 38894
rect 49756 38834 49812 39116
rect 49756 38782 49758 38834
rect 49810 38782 49812 38834
rect 49756 38770 49812 38782
rect 50764 38724 50820 38734
rect 50876 38724 50932 39678
rect 52780 39732 52836 42028
rect 53452 41300 53508 42588
rect 53676 42644 53732 43596
rect 53564 42530 53620 42542
rect 53564 42478 53566 42530
rect 53618 42478 53620 42530
rect 53676 42512 53732 42588
rect 53564 41748 53620 42478
rect 53788 42084 53844 44158
rect 54460 44212 54516 45052
rect 55020 44434 55076 45948
rect 55244 45218 55300 46620
rect 55468 46610 55524 46620
rect 56028 46450 56084 46462
rect 56028 46398 56030 46450
rect 56082 46398 56084 46450
rect 56028 46114 56084 46398
rect 56028 46062 56030 46114
rect 56082 46062 56084 46114
rect 55916 46004 55972 46014
rect 56028 46004 56084 46062
rect 55916 46002 56084 46004
rect 55916 45950 55918 46002
rect 55970 45950 56084 46002
rect 55916 45948 56084 45950
rect 55916 45938 55972 45948
rect 55244 45166 55246 45218
rect 55298 45166 55300 45218
rect 55244 45154 55300 45166
rect 55580 45666 55636 45678
rect 55580 45614 55582 45666
rect 55634 45614 55636 45666
rect 55580 45108 55636 45614
rect 55804 45108 55860 45118
rect 55580 45106 55860 45108
rect 55580 45054 55806 45106
rect 55858 45054 55860 45106
rect 55580 45052 55860 45054
rect 55020 44382 55022 44434
rect 55074 44382 55076 44434
rect 55020 44370 55076 44382
rect 54460 44146 54516 44156
rect 54684 42868 54740 42878
rect 54236 42644 54292 42654
rect 54236 42550 54292 42588
rect 54348 42532 54404 42542
rect 54236 42084 54292 42094
rect 53788 42082 54292 42084
rect 53788 42030 54238 42082
rect 54290 42030 54292 42082
rect 53788 42028 54292 42030
rect 54236 42018 54292 42028
rect 53676 41972 53732 41982
rect 53676 41878 53732 41916
rect 54348 41970 54404 42476
rect 54348 41918 54350 41970
rect 54402 41918 54404 41970
rect 54348 41906 54404 41918
rect 53900 41860 53956 41870
rect 53900 41766 53956 41804
rect 54124 41860 54180 41870
rect 54124 41766 54180 41804
rect 53564 41682 53620 41692
rect 54572 41746 54628 41758
rect 54572 41694 54574 41746
rect 54626 41694 54628 41746
rect 54572 41412 54628 41694
rect 54572 41346 54628 41356
rect 53900 41300 53956 41310
rect 53452 41298 53956 41300
rect 53452 41246 53454 41298
rect 53506 41246 53902 41298
rect 53954 41246 53956 41298
rect 53452 41244 53956 41246
rect 53452 41234 53508 41244
rect 53900 41234 53956 41244
rect 54684 41298 54740 42812
rect 55244 42642 55300 42654
rect 55244 42590 55246 42642
rect 55298 42590 55300 42642
rect 55244 42532 55300 42590
rect 54796 41748 54852 41758
rect 54796 41654 54852 41692
rect 54684 41246 54686 41298
rect 54738 41246 54740 41298
rect 54684 41234 54740 41246
rect 55132 41298 55188 41310
rect 55132 41246 55134 41298
rect 55186 41246 55188 41298
rect 52780 39666 52836 39676
rect 53452 40404 53508 40414
rect 50764 38722 50932 38724
rect 50764 38670 50766 38722
rect 50818 38670 50932 38722
rect 50764 38668 50932 38670
rect 52892 38724 52948 38734
rect 50764 38658 50820 38668
rect 52892 38630 52948 38668
rect 53452 38162 53508 40348
rect 55132 40402 55188 41246
rect 55132 40350 55134 40402
rect 55186 40350 55188 40402
rect 55132 40338 55188 40350
rect 53676 38836 53732 38846
rect 53676 38742 53732 38780
rect 54572 38836 54628 38846
rect 54236 38724 54292 38734
rect 54236 38630 54292 38668
rect 54572 38722 54628 38780
rect 55244 38836 55300 42476
rect 55804 42532 55860 45052
rect 56140 42868 56196 48860
rect 56252 47684 56308 49644
rect 56588 49634 56644 49644
rect 57372 48468 57428 48478
rect 57372 48374 57428 48412
rect 56252 46898 56308 47628
rect 56364 48130 56420 48142
rect 56364 48078 56366 48130
rect 56418 48078 56420 48130
rect 56364 47572 56420 48078
rect 56364 47506 56420 47516
rect 57260 47572 57316 47582
rect 57260 47478 57316 47516
rect 57932 47460 57988 49980
rect 58044 49970 58100 49980
rect 58044 49140 58100 49150
rect 58044 49046 58100 49084
rect 58044 48354 58100 48366
rect 58044 48302 58046 48354
rect 58098 48302 58100 48354
rect 58044 47908 58100 48302
rect 58044 47842 58100 47852
rect 56252 46846 56254 46898
rect 56306 46846 56308 46898
rect 56252 46834 56308 46846
rect 57372 47458 57988 47460
rect 57372 47406 57934 47458
rect 57986 47406 57988 47458
rect 57372 47404 57988 47406
rect 56700 46562 56756 46574
rect 56700 46510 56702 46562
rect 56754 46510 56756 46562
rect 56700 46450 56756 46510
rect 56700 46398 56702 46450
rect 56754 46398 56756 46450
rect 56700 46386 56756 46398
rect 57260 46452 57316 46462
rect 57260 45444 57316 46396
rect 57372 46004 57428 47404
rect 57932 47394 57988 47404
rect 57484 46900 57540 46910
rect 57484 46806 57540 46844
rect 58044 46786 58100 46798
rect 58044 46734 58046 46786
rect 58098 46734 58100 46786
rect 58044 46564 58100 46734
rect 58044 46498 58100 46508
rect 57372 46002 57540 46004
rect 57372 45950 57374 46002
rect 57426 45950 57540 46002
rect 57372 45948 57540 45950
rect 57372 45938 57428 45948
rect 57260 45388 57428 45444
rect 56364 45108 56420 45118
rect 56252 45052 56364 45108
rect 56252 43652 56308 45052
rect 56364 45014 56420 45052
rect 57260 44210 57316 44222
rect 57260 44158 57262 44210
rect 57314 44158 57316 44210
rect 57260 43708 57316 44158
rect 56252 42980 56308 43596
rect 56252 42914 56308 42924
rect 57148 43652 57316 43708
rect 57148 43316 57204 43652
rect 57260 43316 57316 43326
rect 57148 43314 57316 43316
rect 57148 43262 57262 43314
rect 57314 43262 57316 43314
rect 57148 43260 57316 43262
rect 56140 42802 56196 42812
rect 56364 42868 56420 42878
rect 56364 42774 56420 42812
rect 55804 42466 55860 42476
rect 56812 42532 56868 42542
rect 56812 42438 56868 42476
rect 56028 40964 56084 40974
rect 56028 40514 56084 40908
rect 56028 40462 56030 40514
rect 56082 40462 56084 40514
rect 56028 40450 56084 40462
rect 55244 38770 55300 38780
rect 54572 38670 54574 38722
rect 54626 38670 54628 38722
rect 53452 38110 53454 38162
rect 53506 38110 53508 38162
rect 53452 38098 53508 38110
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 53564 37492 53620 37502
rect 53564 37398 53620 37436
rect 54012 37492 54068 37502
rect 54012 37378 54068 37436
rect 54012 37326 54014 37378
rect 54066 37326 54068 37378
rect 54012 37314 54068 37326
rect 54348 37378 54404 37390
rect 54348 37326 54350 37378
rect 54402 37326 54404 37378
rect 49532 37202 49588 37212
rect 48300 36542 48302 36594
rect 48354 36542 48356 36594
rect 48300 36530 48356 36542
rect 50428 36594 50484 36606
rect 50428 36542 50430 36594
rect 50482 36542 50484 36594
rect 42812 26462 42814 26514
rect 42866 26462 42868 26514
rect 42252 26404 42308 26414
rect 42252 26402 42644 26404
rect 42252 26350 42254 26402
rect 42306 26350 42644 26402
rect 42252 26348 42644 26350
rect 42252 26338 42308 26348
rect 42028 26292 42084 26302
rect 42028 26198 42084 26236
rect 42588 25618 42644 26348
rect 42812 26292 42868 26462
rect 42812 26226 42868 26236
rect 47516 36484 47572 36494
rect 42588 25566 42590 25618
rect 42642 25566 42644 25618
rect 42588 25554 42644 25566
rect 43932 25620 43988 25630
rect 43372 25506 43428 25518
rect 43372 25454 43374 25506
rect 43426 25454 43428 25506
rect 43372 25284 43428 25454
rect 43372 25218 43428 25228
rect 43932 25284 43988 25564
rect 47516 25620 47572 36428
rect 47516 25554 47572 25564
rect 43932 25218 43988 25228
rect 50428 4564 50484 36542
rect 50876 36484 50932 36494
rect 50876 36390 50932 36428
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 54348 35812 54404 37326
rect 54348 35746 54404 35756
rect 54572 36484 54628 38670
rect 54572 35364 54628 36428
rect 54572 35026 54628 35308
rect 54572 34974 54574 35026
rect 54626 34974 54628 35026
rect 54572 34962 54628 34974
rect 54796 38724 54852 38734
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 54796 20188 54852 38668
rect 56364 38050 56420 38062
rect 56364 37998 56366 38050
rect 56418 37998 56420 38050
rect 55580 37938 55636 37950
rect 55580 37886 55582 37938
rect 55634 37886 55636 37938
rect 55132 37156 55188 37166
rect 55580 37156 55636 37886
rect 56364 37828 56420 37998
rect 56812 37828 56868 37838
rect 56364 37826 56868 37828
rect 56364 37774 56814 37826
rect 56866 37774 56868 37826
rect 56364 37772 56868 37774
rect 55132 37154 55636 37156
rect 55132 37102 55134 37154
rect 55186 37102 55636 37154
rect 55132 37100 55636 37102
rect 56252 37378 56308 37390
rect 56252 37326 56254 37378
rect 56306 37326 56308 37378
rect 56252 37156 56308 37326
rect 55132 37090 55188 37100
rect 56252 37090 56308 37100
rect 54908 36484 54964 36494
rect 54908 36370 54964 36428
rect 56364 36484 56420 37772
rect 56812 37762 56868 37772
rect 56364 36418 56420 36428
rect 54908 36318 54910 36370
rect 54962 36318 54964 36370
rect 54908 36306 54964 36318
rect 55244 36260 55300 36270
rect 55132 35364 55188 35374
rect 55132 34914 55188 35308
rect 55132 34862 55134 34914
rect 55186 34862 55188 34914
rect 55132 34850 55188 34862
rect 55132 23156 55188 23166
rect 55132 23042 55188 23100
rect 55132 22990 55134 23042
rect 55186 22990 55188 23042
rect 55132 22978 55188 22990
rect 54796 20132 54964 20188
rect 54908 19906 54964 20132
rect 54908 19854 54910 19906
rect 54962 19854 54964 19906
rect 54908 19842 54964 19854
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 55244 8428 55300 36204
rect 55804 36260 55860 36270
rect 55804 36166 55860 36204
rect 55916 35812 55972 35822
rect 55356 35586 55412 35598
rect 55356 35534 55358 35586
rect 55410 35534 55412 35586
rect 55356 35140 55412 35534
rect 55356 35074 55412 35084
rect 55916 35026 55972 35756
rect 55916 34974 55918 35026
rect 55970 34974 55972 35026
rect 55916 34962 55972 34974
rect 56140 35698 56196 35710
rect 56140 35646 56142 35698
rect 56194 35646 56196 35698
rect 56140 35028 56196 35646
rect 56140 34962 56196 34972
rect 56252 23266 56308 23278
rect 56252 23214 56254 23266
rect 56306 23214 56308 23266
rect 56252 23044 56308 23214
rect 57148 23156 57204 43260
rect 57260 43250 57316 43260
rect 57260 41300 57316 41310
rect 57372 41300 57428 45388
rect 57484 45108 57540 45948
rect 58044 45668 58100 45678
rect 58044 45574 58100 45612
rect 57484 45042 57540 45052
rect 58044 45218 58100 45230
rect 58044 45166 58046 45218
rect 58098 45166 58100 45218
rect 58044 44548 58100 45166
rect 58044 44482 58100 44492
rect 57932 44322 57988 44334
rect 57932 44270 57934 44322
rect 57986 44270 57988 44322
rect 57596 43652 57652 43662
rect 57596 43558 57652 43596
rect 57932 43652 57988 44270
rect 57932 43586 57988 43596
rect 58044 43426 58100 43438
rect 58044 43374 58046 43426
rect 58098 43374 58100 43426
rect 58044 43314 58100 43374
rect 58044 43262 58046 43314
rect 58098 43262 58100 43314
rect 58044 43250 58100 43262
rect 57260 41298 57428 41300
rect 57260 41246 57262 41298
rect 57314 41246 57428 41298
rect 57260 41244 57428 41246
rect 57932 42868 57988 42878
rect 57260 41234 57316 41244
rect 57932 41186 57988 42812
rect 57932 41134 57934 41186
rect 57986 41134 57988 41186
rect 57932 41122 57988 41134
rect 58044 40516 58100 40526
rect 58044 40422 58100 40460
rect 58044 39394 58100 39406
rect 58044 39342 58046 39394
rect 58098 39342 58100 39394
rect 58044 39172 58100 39342
rect 58044 39106 58100 39116
rect 57372 37156 57428 37166
rect 57372 37062 57428 37100
rect 58044 35028 58100 35038
rect 58044 34934 58100 34972
rect 57372 31554 57428 31566
rect 57372 31502 57374 31554
rect 57426 31502 57428 31554
rect 57372 31108 57428 31502
rect 58044 31556 58100 31566
rect 58044 31462 58100 31500
rect 57372 31042 57428 31052
rect 58044 31106 58100 31118
rect 58044 31054 58046 31106
rect 58098 31054 58100 31106
rect 58044 30436 58100 31054
rect 58044 30370 58100 30380
rect 58044 28420 58100 28430
rect 58044 28326 58100 28364
rect 58044 24834 58100 24846
rect 58044 24782 58046 24834
rect 58098 24782 58100 24834
rect 58044 24388 58100 24782
rect 58044 24322 58100 24332
rect 57148 23090 57204 23100
rect 56252 22978 56308 22988
rect 57372 23044 57428 23054
rect 57372 22950 57428 22988
rect 56252 20130 56308 20142
rect 56252 20078 56254 20130
rect 56306 20078 56308 20130
rect 56252 19684 56308 20078
rect 56252 19618 56308 19628
rect 57372 19906 57428 19918
rect 57372 19854 57374 19906
rect 57426 19854 57428 19906
rect 57372 19684 57428 19854
rect 57372 19618 57428 19628
rect 58044 15874 58100 15886
rect 58044 15822 58046 15874
rect 58098 15822 58100 15874
rect 58044 15652 58100 15822
rect 58044 15586 58100 15596
rect 58044 13858 58100 13870
rect 58044 13806 58046 13858
rect 58098 13806 58100 13858
rect 58044 13636 58100 13806
rect 58044 13570 58100 13580
rect 58044 11170 58100 11182
rect 58044 11118 58046 11170
rect 58098 11118 58100 11170
rect 58044 10948 58100 11118
rect 58044 10882 58100 10892
rect 55132 8372 55300 8428
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50764 4564 50820 4574
rect 50428 4562 50820 4564
rect 50428 4510 50766 4562
rect 50818 4510 50820 4562
rect 50428 4508 50820 4510
rect 40908 3602 40964 3612
rect 50540 3554 50596 4508
rect 50764 4498 50820 4508
rect 55132 4226 55188 8372
rect 58044 6018 58100 6030
rect 58044 5966 58046 6018
rect 58098 5966 58100 6018
rect 58044 5572 58100 5966
rect 58044 5506 58100 5516
rect 58044 4900 58100 4910
rect 58044 4898 58212 4900
rect 58044 4846 58046 4898
rect 58098 4846 58212 4898
rect 58044 4844 58212 4846
rect 58044 4834 58100 4844
rect 55132 4174 55134 4226
rect 55186 4174 55188 4226
rect 55132 4162 55188 4174
rect 56252 4450 56308 4462
rect 56252 4398 56254 4450
rect 56306 4398 56308 4450
rect 56252 4228 56308 4398
rect 58044 4450 58100 4462
rect 58044 4398 58046 4450
rect 58098 4398 58100 4450
rect 56252 4162 56308 4172
rect 57372 4228 57428 4238
rect 57372 4134 57428 4172
rect 50540 3502 50542 3554
rect 50594 3502 50596 3554
rect 50540 3490 50596 3502
rect 58044 3556 58100 4398
rect 58044 3490 58100 3500
rect 28588 3444 28644 3454
rect 28476 3388 28588 3444
rect 12908 3332 12964 3342
rect 12908 800 12964 3276
rect 13580 3332 13636 3342
rect 15036 3332 15092 3342
rect 16380 3332 16436 3342
rect 19068 3332 19124 3342
rect 22428 3332 22484 3342
rect 23100 3332 23156 3342
rect 24444 3332 24500 3342
rect 28476 3332 28532 3388
rect 13580 3238 13636 3276
rect 14924 3330 15092 3332
rect 14924 3278 15038 3330
rect 15090 3278 15092 3330
rect 14924 3276 15092 3278
rect 14924 800 14980 3276
rect 15036 3266 15092 3276
rect 16268 3330 16436 3332
rect 16268 3278 16382 3330
rect 16434 3278 16436 3330
rect 16268 3276 16436 3278
rect 16268 800 16324 3276
rect 16380 3266 16436 3276
rect 18956 3330 19124 3332
rect 18956 3278 19070 3330
rect 19122 3278 19124 3330
rect 18956 3276 19124 3278
rect 18956 800 19012 3276
rect 19068 3266 19124 3276
rect 22316 3330 22484 3332
rect 22316 3278 22430 3330
rect 22482 3278 22484 3330
rect 22316 3276 22484 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22316 800 22372 3276
rect 22428 3266 22484 3276
rect 22988 3330 23156 3332
rect 22988 3278 23102 3330
rect 23154 3278 23156 3330
rect 22988 3276 23156 3278
rect 22988 800 23044 3276
rect 23100 3266 23156 3276
rect 24332 3330 24500 3332
rect 24332 3278 24446 3330
rect 24498 3278 24500 3330
rect 24332 3276 24500 3278
rect 24332 800 24388 3276
rect 24444 3266 24500 3276
rect 28364 3276 28532 3332
rect 28588 3312 28644 3388
rect 29372 3444 29428 3454
rect 49420 3444 49476 3454
rect 29372 3350 29428 3388
rect 49196 3442 49476 3444
rect 49196 3390 49422 3442
rect 49474 3390 49476 3442
rect 49196 3388 49476 3390
rect 33180 3330 33236 3342
rect 35196 3332 35252 3342
rect 33180 3278 33182 3330
rect 33234 3278 33236 3330
rect 28364 800 28420 3276
rect 32396 1762 32452 1774
rect 32396 1710 32398 1762
rect 32450 1710 32452 1762
rect 32396 800 32452 1710
rect 33180 1762 33236 3278
rect 33180 1710 33182 1762
rect 33234 1710 33236 1762
rect 33180 1698 33236 1710
rect 35084 3330 35252 3332
rect 35084 3278 35198 3330
rect 35250 3278 35252 3330
rect 35084 3276 35252 3278
rect 35084 800 35140 3276
rect 35196 3266 35252 3276
rect 36428 3332 36484 3342
rect 36428 800 36484 3276
rect 37100 3332 37156 3342
rect 39228 3332 39284 3342
rect 39900 3332 39956 3342
rect 46620 3332 46676 3342
rect 47292 3332 47348 3342
rect 37100 3238 37156 3276
rect 39116 3330 39284 3332
rect 39116 3278 39230 3330
rect 39282 3278 39284 3330
rect 39116 3276 39284 3278
rect 39116 800 39172 3276
rect 39228 3266 39284 3276
rect 39788 3330 39956 3332
rect 39788 3278 39902 3330
rect 39954 3278 39956 3330
rect 39788 3276 39956 3278
rect 39788 800 39844 3276
rect 39900 3266 39956 3276
rect 46508 3330 46676 3332
rect 46508 3278 46622 3330
rect 46674 3278 46676 3330
rect 46508 3276 46676 3278
rect 46508 800 46564 3276
rect 46620 3266 46676 3276
rect 47180 3330 47348 3332
rect 47180 3278 47294 3330
rect 47346 3278 47348 3330
rect 47180 3276 47348 3278
rect 47180 800 47236 3276
rect 47292 3266 47348 3276
rect 48076 3332 48132 3342
rect 48076 3330 48356 3332
rect 48076 3278 48078 3330
rect 48130 3278 48356 3330
rect 48076 3276 48356 3278
rect 48076 3266 48132 3276
rect 48300 800 48356 3276
rect 49196 800 49252 3388
rect 49420 3378 49476 3388
rect 51100 3330 51156 3342
rect 51100 3278 51102 3330
rect 51154 3278 51156 3330
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50540 1762 50596 1774
rect 50540 1710 50542 1762
rect 50594 1710 50596 1762
rect 50540 800 50596 1710
rect 51100 1762 51156 3278
rect 51100 1710 51102 1762
rect 51154 1710 51156 1762
rect 51100 1698 51156 1710
rect 51772 3330 51828 3342
rect 51772 3278 51774 3330
rect 51826 3278 51828 3330
rect 51212 812 51380 868
rect 51212 800 51268 812
rect -56 728 196 800
rect -56 200 168 728
rect 616 200 840 800
rect 1288 728 1540 800
rect 1288 200 1512 728
rect 1960 200 2184 800
rect 2632 200 2856 800
rect 3304 728 3556 800
rect 3976 728 4228 800
rect 3304 200 3528 728
rect 3976 200 4200 728
rect 4648 200 4872 800
rect 5320 200 5544 800
rect 5992 200 6216 800
rect 6664 200 6888 800
rect 7336 200 7560 800
rect 8680 200 8904 800
rect 9352 200 9576 800
rect 10024 200 10248 800
rect 10696 200 10920 800
rect 11368 728 11620 800
rect 12040 728 12292 800
rect 12712 728 12964 800
rect 11368 200 11592 728
rect 12040 200 12264 728
rect 12712 200 12936 728
rect 13384 200 13608 800
rect 14056 200 14280 800
rect 14728 728 14980 800
rect 14728 200 14952 728
rect 15400 200 15624 800
rect 16072 728 16324 800
rect 16072 200 16296 728
rect 17416 200 17640 800
rect 18088 200 18312 800
rect 18760 728 19012 800
rect 18760 200 18984 728
rect 19432 200 19656 800
rect 20104 200 20328 800
rect 20776 200 21000 800
rect 21448 200 21672 800
rect 22120 728 22372 800
rect 22792 728 23044 800
rect 22120 200 22344 728
rect 22792 200 23016 728
rect 23464 200 23688 800
rect 24136 728 24388 800
rect 24136 200 24360 728
rect 24808 200 25032 800
rect 26152 200 26376 800
rect 26824 200 27048 800
rect 27496 200 27720 800
rect 28168 728 28420 800
rect 28168 200 28392 728
rect 28840 200 29064 800
rect 29512 200 29736 800
rect 30184 200 30408 800
rect 30856 200 31080 800
rect 31528 200 31752 800
rect 32200 728 32452 800
rect 32200 200 32424 728
rect 32872 200 33096 800
rect 33544 200 33768 800
rect 34888 728 35140 800
rect 34888 200 35112 728
rect 35560 200 35784 800
rect 36232 728 36484 800
rect 36232 200 36456 728
rect 36904 200 37128 800
rect 37576 200 37800 800
rect 38248 200 38472 800
rect 38920 728 39172 800
rect 39592 728 39844 800
rect 38920 200 39144 728
rect 39592 200 39816 728
rect 40264 200 40488 800
rect 40936 200 41160 800
rect 41608 200 41832 800
rect 42280 200 42504 800
rect 43624 200 43848 800
rect 44296 200 44520 800
rect 44968 200 45192 800
rect 45640 200 45864 800
rect 46312 728 46564 800
rect 46984 728 47236 800
rect 46312 200 46536 728
rect 46984 200 47208 728
rect 47656 200 47880 800
rect 48300 728 48552 800
rect 48328 200 48552 728
rect 49000 728 49252 800
rect 49000 200 49224 728
rect 49672 200 49896 800
rect 50344 728 50596 800
rect 51016 728 51268 800
rect 51324 756 51380 812
rect 51772 756 51828 3278
rect 55916 3330 55972 3342
rect 55916 3278 55918 3330
rect 55970 3278 55972 3330
rect 55916 2212 55972 3278
rect 55916 2146 55972 2156
rect 56700 3330 56756 3342
rect 56700 3278 56702 3330
rect 56754 3278 56756 3330
rect 55916 1762 55972 1774
rect 55916 1710 55918 1762
rect 55970 1710 55972 1762
rect 55916 800 55972 1710
rect 56700 1762 56756 3278
rect 56700 1710 56702 1762
rect 56754 1710 56756 1762
rect 56700 1698 56756 1710
rect 57932 3330 57988 3342
rect 57932 3278 57934 3330
rect 57986 3278 57988 3330
rect 57932 800 57988 3278
rect 50344 200 50568 728
rect 51016 200 51240 728
rect 51324 700 51828 756
rect 52360 200 52584 800
rect 53032 200 53256 800
rect 53704 200 53928 800
rect 54376 200 54600 800
rect 55048 200 55272 800
rect 55720 728 55972 800
rect 55720 200 55944 728
rect 56392 200 56616 800
rect 57064 200 57288 800
rect 57736 728 57988 800
rect 57736 200 57960 728
rect 58156 196 58212 4844
rect 58408 200 58632 800
rect 59080 200 59304 800
rect 58156 130 58212 140
<< via2 >>
rect 3164 58380 3220 58436
rect 1820 55244 1876 55300
rect 3052 55298 3108 55300
rect 3052 55246 3054 55298
rect 3054 55246 3106 55298
rect 3106 55246 3108 55298
rect 3052 55244 3108 55246
rect 1484 54684 1540 54740
rect 2492 54738 2548 54740
rect 2492 54686 2494 54738
rect 2494 54686 2546 54738
rect 2546 54686 2548 54738
rect 2492 54684 2548 54686
rect 4060 57148 4116 57204
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 3724 55244 3780 55300
rect 1932 54572 1988 54628
rect 1820 53900 1876 53956
rect 1932 53228 1988 53284
rect 1820 52556 1876 52612
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 3724 52780 3780 52836
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 3500 51996 3556 52052
rect 1820 51212 1876 51268
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 12796 56082 12852 56084
rect 12796 56030 12798 56082
rect 12798 56030 12850 56082
rect 12850 56030 12852 56082
rect 12796 56028 12852 56030
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 36428 56252 36484 56308
rect 37100 56306 37156 56308
rect 37100 56254 37102 56306
rect 37102 56254 37154 56306
rect 37154 56254 37156 56306
rect 37100 56252 37156 56254
rect 46508 56252 46564 56308
rect 47964 56306 48020 56308
rect 47964 56254 47966 56306
rect 47966 56254 48018 56306
rect 48018 56254 48020 56306
rect 47964 56252 48020 56254
rect 57484 58380 57540 58436
rect 56588 56588 56644 56644
rect 57372 56588 57428 56644
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 15036 56082 15092 56084
rect 15036 56030 15038 56082
rect 15038 56030 15090 56082
rect 15090 56030 15092 56082
rect 15036 56028 15092 56030
rect 12908 55132 12964 55188
rect 13692 55186 13748 55188
rect 13692 55134 13694 55186
rect 13694 55134 13746 55186
rect 13746 55134 13748 55186
rect 13692 55132 13748 55134
rect 46284 55916 46340 55972
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 47180 55970 47236 55972
rect 47180 55918 47182 55970
rect 47182 55918 47234 55970
rect 47234 55918 47236 55970
rect 47180 55916 47236 55918
rect 55916 55970 55972 55972
rect 55916 55918 55918 55970
rect 55918 55918 55970 55970
rect 55970 55918 55972 55970
rect 55916 55916 55972 55918
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 15036 54348 15092 54404
rect 41580 54402 41636 54404
rect 41580 54350 41582 54402
rect 41582 54350 41634 54402
rect 41634 54350 41636 54402
rect 41580 54348 41636 54350
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 7196 53452 7252 53508
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 44156 53116 44212 53172
rect 44492 54348 44548 54404
rect 44380 53170 44436 53172
rect 44380 53118 44382 53170
rect 44382 53118 44434 53170
rect 44434 53118 44436 53170
rect 44380 53116 44436 53118
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 42812 52220 42868 52276
rect 39900 51996 39956 52052
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 43260 52274 43316 52276
rect 43260 52222 43262 52274
rect 43262 52222 43314 52274
rect 43314 52222 43316 52274
rect 43260 52220 43316 52222
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 41692 50988 41748 51044
rect 35404 50932 35460 50934
rect 4844 50652 4900 50708
rect 44044 51938 44100 51940
rect 44044 51886 44046 51938
rect 44046 51886 44098 51938
rect 44098 51886 44100 51938
rect 44044 51884 44100 51886
rect 44044 51490 44100 51492
rect 44044 51438 44046 51490
rect 44046 51438 44098 51490
rect 44098 51438 44100 51490
rect 44044 51436 44100 51438
rect 39564 50706 39620 50708
rect 39564 50654 39566 50706
rect 39566 50654 39618 50706
rect 39618 50654 39620 50706
rect 39564 50652 39620 50654
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 44940 54402 44996 54404
rect 44940 54350 44942 54402
rect 44942 54350 44994 54402
rect 44994 54350 44996 54402
rect 44940 54348 44996 54350
rect 45612 54348 45668 54404
rect 45612 53788 45668 53844
rect 47292 53788 47348 53844
rect 44716 53730 44772 53732
rect 44716 53678 44718 53730
rect 44718 53678 44770 53730
rect 44770 53678 44772 53730
rect 44716 53676 44772 53678
rect 47292 53564 47348 53620
rect 46732 53506 46788 53508
rect 46732 53454 46734 53506
rect 46734 53454 46786 53506
rect 46786 53454 46788 53506
rect 46732 53452 46788 53454
rect 47964 53452 48020 53508
rect 45276 53170 45332 53172
rect 45276 53118 45278 53170
rect 45278 53118 45330 53170
rect 45330 53118 45332 53170
rect 45276 53116 45332 53118
rect 44828 53004 44884 53060
rect 44716 52946 44772 52948
rect 44716 52894 44718 52946
rect 44718 52894 44770 52946
rect 44770 52894 44772 52946
rect 44716 52892 44772 52894
rect 44492 52220 44548 52276
rect 45500 53058 45556 53060
rect 45500 53006 45502 53058
rect 45502 53006 45554 53058
rect 45554 53006 45556 53058
rect 45500 53004 45556 53006
rect 48076 53058 48132 53060
rect 48076 53006 48078 53058
rect 48078 53006 48130 53058
rect 48130 53006 48132 53058
rect 48076 53004 48132 53006
rect 45612 52946 45668 52948
rect 45612 52894 45614 52946
rect 45614 52894 45666 52946
rect 45666 52894 45668 52946
rect 45612 52892 45668 52894
rect 44604 51324 44660 51380
rect 44716 51884 44772 51940
rect 44828 51772 44884 51828
rect 44828 51490 44884 51492
rect 44828 51438 44830 51490
rect 44830 51438 44882 51490
rect 44882 51438 44884 51490
rect 44828 51436 44884 51438
rect 45724 51938 45780 51940
rect 45724 51886 45726 51938
rect 45726 51886 45778 51938
rect 45778 51886 45780 51938
rect 45724 51884 45780 51886
rect 46732 51996 46788 52052
rect 46396 51938 46452 51940
rect 46396 51886 46398 51938
rect 46398 51886 46450 51938
rect 46450 51886 46452 51938
rect 46396 51884 46452 51886
rect 46396 51660 46452 51716
rect 45836 51490 45892 51492
rect 45836 51438 45838 51490
rect 45838 51438 45890 51490
rect 45890 51438 45892 51490
rect 45836 51436 45892 51438
rect 45948 51378 46004 51380
rect 45948 51326 45950 51378
rect 45950 51326 46002 51378
rect 46002 51326 46004 51378
rect 45948 51324 46004 51326
rect 46396 51378 46452 51380
rect 46396 51326 46398 51378
rect 46398 51326 46450 51378
rect 46450 51326 46452 51378
rect 46396 51324 46452 51326
rect 46284 50706 46340 50708
rect 46284 50654 46286 50706
rect 46286 50654 46338 50706
rect 46338 50654 46340 50706
rect 46284 50652 46340 50654
rect 45388 50540 45444 50596
rect 44716 50482 44772 50484
rect 44716 50430 44718 50482
rect 44718 50430 44770 50482
rect 44770 50430 44772 50482
rect 44716 50428 44772 50430
rect 47292 52050 47348 52052
rect 47292 51998 47294 52050
rect 47294 51998 47346 52050
rect 47346 51998 47348 52050
rect 47292 51996 47348 51998
rect 46732 50652 46788 50708
rect 45276 50428 45332 50484
rect 44268 49756 44324 49812
rect 42700 49138 42756 49140
rect 42700 49086 42702 49138
rect 42702 49086 42754 49138
rect 42754 49086 42756 49138
rect 42700 49084 42756 49086
rect 44604 49810 44660 49812
rect 44604 49758 44606 49810
rect 44606 49758 44658 49810
rect 44658 49758 44660 49810
rect 44604 49756 44660 49758
rect 44940 49810 44996 49812
rect 44940 49758 44942 49810
rect 44942 49758 44994 49810
rect 44994 49758 44996 49810
rect 44940 49756 44996 49758
rect 44268 49084 44324 49140
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 44156 48860 44212 48916
rect 44492 49026 44548 49028
rect 44492 48974 44494 49026
rect 44494 48974 44546 49026
rect 44546 48974 44548 49026
rect 44492 48972 44548 48974
rect 43260 47628 43316 47684
rect 44268 47682 44324 47684
rect 44268 47630 44270 47682
rect 44270 47630 44322 47682
rect 44322 47630 44324 47682
rect 44268 47628 44324 47630
rect 43148 47570 43204 47572
rect 43148 47518 43150 47570
rect 43150 47518 43202 47570
rect 43202 47518 43204 47570
rect 43148 47516 43204 47518
rect 44380 47516 44436 47572
rect 1820 47234 1876 47236
rect 1820 47182 1822 47234
rect 1822 47182 1874 47234
rect 1874 47182 1876 47234
rect 1820 47180 1876 47182
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 43372 47180 43428 47236
rect 44268 47234 44324 47236
rect 44268 47182 44270 47234
rect 44270 47182 44322 47234
rect 44322 47182 44324 47234
rect 44268 47180 44324 47182
rect 43036 46620 43092 46676
rect 42700 45724 42756 45780
rect 2492 45666 2548 45668
rect 2492 45614 2494 45666
rect 2494 45614 2546 45666
rect 2546 45614 2548 45666
rect 2492 45612 2548 45614
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 1708 45164 1764 45220
rect 42812 45164 42868 45220
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 1820 44492 1876 44548
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 40124 42754 40180 42756
rect 40124 42702 40126 42754
rect 40126 42702 40178 42754
rect 40178 42702 40180 42754
rect 40124 42700 40180 42702
rect 42028 42700 42084 42756
rect 39452 42588 39508 42644
rect 40796 42642 40852 42644
rect 40796 42590 40798 42642
rect 40798 42590 40850 42642
rect 40850 42590 40852 42642
rect 40796 42588 40852 42590
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 2492 40962 2548 40964
rect 2492 40910 2494 40962
rect 2494 40910 2546 40962
rect 2546 40910 2548 40962
rect 2492 40908 2548 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 1708 40460 1764 40516
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 1820 39788 1876 39844
rect 1820 39116 1876 39172
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 1820 35084 1876 35140
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 1820 31554 1876 31556
rect 1820 31502 1822 31554
rect 1822 31502 1874 31554
rect 1874 31502 1876 31554
rect 1820 31500 1876 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 2492 31052 2548 31108
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 1820 28418 1876 28420
rect 1820 28366 1822 28418
rect 1822 28366 1874 28418
rect 1874 28366 1876 28418
rect 1820 28364 1876 28366
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 1820 26908 1876 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 3052 25228 3108 25284
rect 3612 25282 3668 25284
rect 3612 25230 3614 25282
rect 3614 25230 3666 25282
rect 3666 25230 3668 25282
rect 3612 25228 3668 25230
rect 1932 25004 1988 25060
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 1820 22988 1876 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 1708 21644 1764 21700
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 1820 20972 1876 21028
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 1820 19628 1876 19684
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 1820 18284 1876 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 1820 16268 1876 16324
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 1820 14924 1876 14980
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 1820 14306 1876 14308
rect 1820 14254 1822 14306
rect 1822 14254 1874 14306
rect 1874 14254 1876 14306
rect 1820 14252 1876 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 1820 12738 1876 12740
rect 1820 12686 1822 12738
rect 1822 12686 1874 12738
rect 1874 12686 1876 12738
rect 1820 12684 1876 12686
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 1820 10220 1876 10276
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 1820 9602 1876 9604
rect 1820 9550 1822 9602
rect 1822 9550 1874 9602
rect 1874 9550 1876 9602
rect 1820 9548 1876 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 1820 6188 1876 6244
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 1820 4898 1876 4900
rect 1820 4846 1822 4898
rect 1822 4846 1874 4898
rect 1874 4846 1876 4898
rect 1820 4844 1876 4846
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 140 1596 196 1652
rect 11564 4172 11620 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 1932 2156 1988 2212
rect 2492 1596 2548 1652
rect 13020 4226 13076 4228
rect 13020 4174 13022 4226
rect 13022 4174 13074 4226
rect 13074 4174 13076 4226
rect 13020 4172 13076 4174
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 30716 3724 30772 3780
rect 12796 3666 12852 3668
rect 12796 3614 12798 3666
rect 12798 3614 12850 3666
rect 12850 3614 12852 3666
rect 12796 3612 12852 3614
rect 40908 40402 40964 40404
rect 40908 40350 40910 40402
rect 40910 40350 40962 40402
rect 40962 40350 40964 40402
rect 40908 40348 40964 40350
rect 40460 25228 40516 25284
rect 39452 3724 39508 3780
rect 42364 40402 42420 40404
rect 42364 40350 42366 40402
rect 42366 40350 42418 40402
rect 42418 40350 42420 40402
rect 42364 40348 42420 40350
rect 43148 45778 43204 45780
rect 43148 45726 43150 45778
rect 43150 45726 43202 45778
rect 43202 45726 43204 45778
rect 43148 45724 43204 45726
rect 43596 45218 43652 45220
rect 43596 45166 43598 45218
rect 43598 45166 43650 45218
rect 43650 45166 43652 45218
rect 43596 45164 43652 45166
rect 44268 45106 44324 45108
rect 44268 45054 44270 45106
rect 44270 45054 44322 45106
rect 44322 45054 44324 45106
rect 44268 45052 44324 45054
rect 43708 44380 43764 44436
rect 44492 44940 44548 44996
rect 43484 44210 43540 44212
rect 43484 44158 43486 44210
rect 43486 44158 43538 44210
rect 43538 44158 43540 44210
rect 43484 44156 43540 44158
rect 44716 44828 44772 44884
rect 44604 44322 44660 44324
rect 44604 44270 44606 44322
rect 44606 44270 44658 44322
rect 44658 44270 44660 44322
rect 44604 44268 44660 44270
rect 44044 44044 44100 44100
rect 43596 42754 43652 42756
rect 43596 42702 43598 42754
rect 43598 42702 43650 42754
rect 43650 42702 43652 42754
rect 43596 42700 43652 42702
rect 44492 40572 44548 40628
rect 45052 45052 45108 45108
rect 45052 44044 45108 44100
rect 44940 42924 44996 42980
rect 46396 49980 46452 50036
rect 45612 49810 45668 49812
rect 45612 49758 45614 49810
rect 45614 49758 45666 49810
rect 45666 49758 45668 49810
rect 45612 49756 45668 49758
rect 45500 48972 45556 49028
rect 45836 49026 45892 49028
rect 45836 48974 45838 49026
rect 45838 48974 45890 49026
rect 45890 48974 45892 49026
rect 45836 48972 45892 48974
rect 45948 48914 46004 48916
rect 45948 48862 45950 48914
rect 45950 48862 46002 48914
rect 46002 48862 46004 48914
rect 45948 48860 46004 48862
rect 46508 48972 46564 49028
rect 46396 48524 46452 48580
rect 46396 48188 46452 48244
rect 45500 47570 45556 47572
rect 45500 47518 45502 47570
rect 45502 47518 45554 47570
rect 45554 47518 45556 47570
rect 45500 47516 45556 47518
rect 47292 50428 47348 50484
rect 47404 50034 47460 50036
rect 47404 49982 47406 50034
rect 47406 49982 47458 50034
rect 47458 49982 47460 50034
rect 47404 49980 47460 49982
rect 48188 51884 48244 51940
rect 48300 51548 48356 51604
rect 48188 51436 48244 51492
rect 47964 50428 48020 50484
rect 48188 50988 48244 51044
rect 47964 49810 48020 49812
rect 47964 49758 47966 49810
rect 47966 49758 48018 49810
rect 48018 49758 48020 49810
rect 47964 49756 48020 49758
rect 47180 48972 47236 49028
rect 46956 48914 47012 48916
rect 46956 48862 46958 48914
rect 46958 48862 47010 48914
rect 47010 48862 47012 48914
rect 46956 48860 47012 48862
rect 47180 48748 47236 48804
rect 47068 48300 47124 48356
rect 46732 48242 46788 48244
rect 46732 48190 46734 48242
rect 46734 48190 46786 48242
rect 46786 48190 46788 48242
rect 46732 48188 46788 48190
rect 46172 47458 46228 47460
rect 46172 47406 46174 47458
rect 46174 47406 46226 47458
rect 46226 47406 46228 47458
rect 46172 47404 46228 47406
rect 47068 47404 47124 47460
rect 46396 47180 46452 47236
rect 46172 46786 46228 46788
rect 46172 46734 46174 46786
rect 46174 46734 46226 46786
rect 46226 46734 46228 46786
rect 46172 46732 46228 46734
rect 46060 44994 46116 44996
rect 46060 44942 46062 44994
rect 46062 44942 46114 44994
rect 46114 44942 46116 44994
rect 46060 44940 46116 44942
rect 45500 44434 45556 44436
rect 45500 44382 45502 44434
rect 45502 44382 45554 44434
rect 45554 44382 45556 44434
rect 45500 44380 45556 44382
rect 45836 44882 45892 44884
rect 45836 44830 45838 44882
rect 45838 44830 45890 44882
rect 45890 44830 45892 44882
rect 45836 44828 45892 44830
rect 46732 46732 46788 46788
rect 46508 46674 46564 46676
rect 46508 46622 46510 46674
rect 46510 46622 46562 46674
rect 46562 46622 46564 46674
rect 46508 46620 46564 46622
rect 54012 55356 54068 55412
rect 55020 55356 55076 55412
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 48860 54684 48916 54740
rect 50540 54684 50596 54740
rect 49420 53004 49476 53060
rect 52220 54626 52276 54628
rect 52220 54574 52222 54626
rect 52222 54574 52274 54626
rect 52274 54574 52276 54626
rect 52220 54572 52276 54574
rect 53564 54626 53620 54628
rect 53564 54574 53566 54626
rect 53566 54574 53618 54626
rect 53618 54574 53620 54626
rect 53564 54572 53620 54574
rect 51884 53676 51940 53732
rect 50540 53618 50596 53620
rect 50540 53566 50542 53618
rect 50542 53566 50594 53618
rect 50594 53566 50596 53618
rect 50540 53564 50596 53566
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 48748 51938 48804 51940
rect 48748 51886 48750 51938
rect 48750 51886 48802 51938
rect 48802 51886 48804 51938
rect 48748 51884 48804 51886
rect 48636 51660 48692 51716
rect 48748 50540 48804 50596
rect 48524 50316 48580 50372
rect 48636 50428 48692 50484
rect 48412 49810 48468 49812
rect 48412 49758 48414 49810
rect 48414 49758 48466 49810
rect 48466 49758 48468 49810
rect 48412 49756 48468 49758
rect 48972 51938 49028 51940
rect 48972 51886 48974 51938
rect 48974 51886 49026 51938
rect 49026 51886 49028 51938
rect 48972 51884 49028 51886
rect 48636 49756 48692 49812
rect 48860 49644 48916 49700
rect 48972 51660 49028 51716
rect 49420 51602 49476 51604
rect 49420 51550 49422 51602
rect 49422 51550 49474 51602
rect 49474 51550 49476 51602
rect 49420 51548 49476 51550
rect 50092 52834 50148 52836
rect 50092 52782 50094 52834
rect 50094 52782 50146 52834
rect 50146 52782 50148 52834
rect 50092 52780 50148 52782
rect 49644 51938 49700 51940
rect 49644 51886 49646 51938
rect 49646 51886 49698 51938
rect 49698 51886 49700 51938
rect 49644 51884 49700 51886
rect 49644 51490 49700 51492
rect 49644 51438 49646 51490
rect 49646 51438 49698 51490
rect 49698 51438 49700 51490
rect 49644 51436 49700 51438
rect 49308 50540 49364 50596
rect 48748 49138 48804 49140
rect 48748 49086 48750 49138
rect 48750 49086 48802 49138
rect 48802 49086 48804 49138
rect 48748 49084 48804 49086
rect 48524 49026 48580 49028
rect 48524 48974 48526 49026
rect 48526 48974 48578 49026
rect 48578 48974 48580 49026
rect 48524 48972 48580 48974
rect 47404 48914 47460 48916
rect 47404 48862 47406 48914
rect 47406 48862 47458 48914
rect 47458 48862 47460 48914
rect 47404 48860 47460 48862
rect 47516 48802 47572 48804
rect 47516 48750 47518 48802
rect 47518 48750 47570 48802
rect 47570 48750 47572 48802
rect 47516 48748 47572 48750
rect 47292 48242 47348 48244
rect 47292 48190 47294 48242
rect 47294 48190 47346 48242
rect 47346 48190 47348 48242
rect 47292 48188 47348 48190
rect 47628 48524 47684 48580
rect 47516 48354 47572 48356
rect 47516 48302 47518 48354
rect 47518 48302 47570 48354
rect 47570 48302 47572 48354
rect 47516 48300 47572 48302
rect 48300 48354 48356 48356
rect 48300 48302 48302 48354
rect 48302 48302 48354 48354
rect 48354 48302 48356 48354
rect 48300 48300 48356 48302
rect 49532 49756 49588 49812
rect 49756 51212 49812 51268
rect 49756 50540 49812 50596
rect 50204 51266 50260 51268
rect 50204 51214 50206 51266
rect 50206 51214 50258 51266
rect 50258 51214 50260 51266
rect 50204 51212 50260 51214
rect 51660 52780 51716 52836
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50652 51436 50708 51492
rect 49644 49868 49700 49924
rect 49084 49532 49140 49588
rect 47068 46786 47124 46788
rect 47068 46734 47070 46786
rect 47070 46734 47122 46786
rect 47122 46734 47124 46786
rect 47068 46732 47124 46734
rect 46956 46620 47012 46676
rect 47292 46674 47348 46676
rect 47292 46622 47294 46674
rect 47294 46622 47346 46674
rect 47346 46622 47348 46674
rect 47292 46620 47348 46622
rect 47516 46396 47572 46452
rect 47068 46284 47124 46340
rect 48300 46956 48356 47012
rect 48188 46898 48244 46900
rect 48188 46846 48190 46898
rect 48190 46846 48242 46898
rect 48242 46846 48244 46898
rect 48188 46844 48244 46846
rect 48748 46956 48804 47012
rect 48524 46674 48580 46676
rect 48524 46622 48526 46674
rect 48526 46622 48578 46674
rect 48578 46622 48580 46674
rect 48524 46620 48580 46622
rect 47628 46284 47684 46340
rect 47068 45724 47124 45780
rect 46732 45388 46788 45444
rect 46508 45106 46564 45108
rect 46508 45054 46510 45106
rect 46510 45054 46562 45106
rect 46562 45054 46564 45106
rect 46508 45052 46564 45054
rect 45948 44322 46004 44324
rect 45948 44270 45950 44322
rect 45950 44270 46002 44322
rect 46002 44270 46004 44322
rect 45948 44268 46004 44270
rect 48188 45890 48244 45892
rect 48188 45838 48190 45890
rect 48190 45838 48242 45890
rect 48242 45838 48244 45890
rect 48188 45836 48244 45838
rect 48860 46620 48916 46676
rect 48748 45948 48804 46004
rect 48412 45778 48468 45780
rect 48412 45726 48414 45778
rect 48414 45726 48466 45778
rect 48466 45726 48468 45778
rect 48412 45724 48468 45726
rect 48636 45612 48692 45668
rect 48188 45106 48244 45108
rect 48188 45054 48190 45106
rect 48190 45054 48242 45106
rect 48242 45054 48244 45106
rect 48188 45052 48244 45054
rect 47964 44940 48020 44996
rect 48972 45388 49028 45444
rect 48524 44828 48580 44884
rect 45388 42812 45444 42868
rect 46284 42866 46340 42868
rect 46284 42814 46286 42866
rect 46286 42814 46338 42866
rect 46338 42814 46340 42866
rect 46284 42812 46340 42814
rect 46172 42530 46228 42532
rect 46172 42478 46174 42530
rect 46174 42478 46226 42530
rect 46226 42478 46228 42530
rect 46172 42476 46228 42478
rect 46396 41970 46452 41972
rect 46396 41918 46398 41970
rect 46398 41918 46450 41970
rect 46450 41918 46452 41970
rect 46396 41916 46452 41918
rect 46620 41356 46676 41412
rect 46732 42476 46788 42532
rect 48748 44156 48804 44212
rect 48972 43372 49028 43428
rect 48524 42866 48580 42868
rect 48524 42814 48526 42866
rect 48526 42814 48578 42866
rect 48578 42814 48580 42866
rect 48524 42812 48580 42814
rect 46620 41186 46676 41188
rect 46620 41134 46622 41186
rect 46622 41134 46674 41186
rect 46674 41134 46676 41186
rect 46620 41132 46676 41134
rect 46396 41020 46452 41076
rect 45276 40572 45332 40628
rect 46284 40626 46340 40628
rect 46284 40574 46286 40626
rect 46286 40574 46338 40626
rect 46338 40574 46340 40626
rect 46284 40572 46340 40574
rect 48076 41916 48132 41972
rect 47964 41692 48020 41748
rect 47404 41410 47460 41412
rect 47404 41358 47406 41410
rect 47406 41358 47458 41410
rect 47458 41358 47460 41410
rect 47404 41356 47460 41358
rect 46844 41132 46900 41188
rect 48076 41356 48132 41412
rect 47292 41186 47348 41188
rect 47292 41134 47294 41186
rect 47294 41134 47346 41186
rect 47346 41134 47348 41186
rect 47292 41132 47348 41134
rect 47404 41074 47460 41076
rect 47404 41022 47406 41074
rect 47406 41022 47458 41074
rect 47458 41022 47460 41074
rect 47404 41020 47460 41022
rect 47068 40572 47124 40628
rect 46956 40514 47012 40516
rect 46956 40462 46958 40514
rect 46958 40462 47010 40514
rect 47010 40462 47012 40514
rect 46956 40460 47012 40462
rect 47404 40460 47460 40516
rect 48300 42530 48356 42532
rect 48300 42478 48302 42530
rect 48302 42478 48354 42530
rect 48354 42478 48356 42530
rect 48300 42476 48356 42478
rect 49980 49644 50036 49700
rect 50652 50428 50708 50484
rect 50876 50370 50932 50372
rect 50876 50318 50878 50370
rect 50878 50318 50930 50370
rect 50930 50318 50932 50370
rect 50876 50316 50932 50318
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50316 49308 50372 49364
rect 50092 49084 50148 49140
rect 49868 48972 49924 49028
rect 49196 48748 49252 48804
rect 49756 48860 49812 48916
rect 49868 48466 49924 48468
rect 49868 48414 49870 48466
rect 49870 48414 49922 48466
rect 49922 48414 49924 48466
rect 49868 48412 49924 48414
rect 49756 47570 49812 47572
rect 49756 47518 49758 47570
rect 49758 47518 49810 47570
rect 49810 47518 49812 47570
rect 49756 47516 49812 47518
rect 49980 47516 50036 47572
rect 49308 46956 49364 47012
rect 49532 46956 49588 47012
rect 49196 45724 49252 45780
rect 49980 46844 50036 46900
rect 50204 48860 50260 48916
rect 50540 48914 50596 48916
rect 50540 48862 50542 48914
rect 50542 48862 50594 48914
rect 50594 48862 50596 48914
rect 50540 48860 50596 48862
rect 50988 49810 51044 49812
rect 50988 49758 50990 49810
rect 50990 49758 51042 49810
rect 51042 49758 51044 49810
rect 50988 49756 51044 49758
rect 52220 52834 52276 52836
rect 52220 52782 52222 52834
rect 52222 52782 52274 52834
rect 52274 52782 52276 52834
rect 52220 52780 52276 52782
rect 56252 55186 56308 55188
rect 56252 55134 56254 55186
rect 56254 55134 56306 55186
rect 56306 55134 56308 55186
rect 56252 55132 56308 55134
rect 56700 55132 56756 55188
rect 55132 52220 55188 52276
rect 55580 52274 55636 52276
rect 55580 52222 55582 52274
rect 55582 52222 55634 52274
rect 55634 52222 55636 52274
rect 55580 52220 55636 52222
rect 57260 55916 57316 55972
rect 52108 50316 52164 50372
rect 51772 49980 51828 50036
rect 51884 50092 51940 50148
rect 51324 49756 51380 49812
rect 51772 49810 51828 49812
rect 51772 49758 51774 49810
rect 51774 49758 51826 49810
rect 51826 49758 51828 49810
rect 51772 49756 51828 49758
rect 51548 49644 51604 49700
rect 51660 49026 51716 49028
rect 51660 48974 51662 49026
rect 51662 48974 51714 49026
rect 51714 48974 51716 49026
rect 51660 48972 51716 48974
rect 50876 48860 50932 48916
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50428 48076 50484 48132
rect 49644 46450 49700 46452
rect 49644 46398 49646 46450
rect 49646 46398 49698 46450
rect 49698 46398 49700 46450
rect 49644 46396 49700 46398
rect 50204 46956 50260 47012
rect 50092 46002 50148 46004
rect 50092 45950 50094 46002
rect 50094 45950 50146 46002
rect 50146 45950 50148 46002
rect 50092 45948 50148 45950
rect 49644 45836 49700 45892
rect 49644 45666 49700 45668
rect 49644 45614 49646 45666
rect 49646 45614 49698 45666
rect 49698 45614 49700 45666
rect 49644 45612 49700 45614
rect 49420 42866 49476 42868
rect 49420 42814 49422 42866
rect 49422 42814 49474 42866
rect 49474 42814 49476 42866
rect 49420 42812 49476 42814
rect 50652 47570 50708 47572
rect 50652 47518 50654 47570
rect 50654 47518 50706 47570
rect 50706 47518 50708 47570
rect 50652 47516 50708 47518
rect 50988 48130 51044 48132
rect 50988 48078 50990 48130
rect 50990 48078 51042 48130
rect 51042 48078 51044 48130
rect 50988 48076 51044 48078
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 51212 47516 51268 47572
rect 50988 46956 51044 47012
rect 51100 46844 51156 46900
rect 50764 46002 50820 46004
rect 50764 45950 50766 46002
rect 50766 45950 50818 46002
rect 50818 45950 50820 46002
rect 50764 45948 50820 45950
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 51548 48524 51604 48580
rect 51996 49308 52052 49364
rect 52556 50092 52612 50148
rect 53004 50204 53060 50260
rect 52668 49196 52724 49252
rect 52220 48972 52276 49028
rect 52556 49026 52612 49028
rect 52556 48974 52558 49026
rect 52558 48974 52610 49026
rect 52610 48974 52612 49026
rect 52556 48972 52612 48974
rect 52108 48412 52164 48468
rect 51436 46956 51492 47012
rect 51548 46898 51604 46900
rect 51548 46846 51550 46898
rect 51550 46846 51602 46898
rect 51602 46846 51604 46898
rect 51548 46844 51604 46846
rect 51324 45836 51380 45892
rect 50988 45612 51044 45668
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 49868 42812 49924 42868
rect 48412 41244 48468 41300
rect 48300 41186 48356 41188
rect 48300 41134 48302 41186
rect 48302 41134 48354 41186
rect 48354 41134 48356 41186
rect 48300 41132 48356 41134
rect 48188 41020 48244 41076
rect 47852 40460 47908 40516
rect 47964 40572 48020 40628
rect 48636 41858 48692 41860
rect 48636 41806 48638 41858
rect 48638 41806 48690 41858
rect 48690 41806 48692 41858
rect 48636 41804 48692 41806
rect 49756 41916 49812 41972
rect 49532 41858 49588 41860
rect 49532 41806 49534 41858
rect 49534 41806 49586 41858
rect 49586 41806 49588 41858
rect 49532 41804 49588 41806
rect 49644 41410 49700 41412
rect 49644 41358 49646 41410
rect 49646 41358 49698 41410
rect 49698 41358 49700 41410
rect 49644 41356 49700 41358
rect 49980 41692 50036 41748
rect 49644 41074 49700 41076
rect 49644 41022 49646 41074
rect 49646 41022 49698 41074
rect 49698 41022 49700 41074
rect 49644 41020 49700 41022
rect 50876 43426 50932 43428
rect 50876 43374 50878 43426
rect 50878 43374 50930 43426
rect 50930 43374 50932 43426
rect 50876 43372 50932 43374
rect 51324 45666 51380 45668
rect 51324 45614 51326 45666
rect 51326 45614 51378 45666
rect 51378 45614 51380 45666
rect 51324 45612 51380 45614
rect 51436 45500 51492 45556
rect 51212 43596 51268 43652
rect 51100 43372 51156 43428
rect 50988 42476 51044 42532
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50428 41916 50484 41972
rect 50316 41692 50372 41748
rect 50876 41692 50932 41748
rect 50204 41020 50260 41076
rect 51996 46620 52052 46676
rect 51884 46396 51940 46452
rect 52780 48636 52836 48692
rect 53004 49922 53060 49924
rect 53004 49870 53006 49922
rect 53006 49870 53058 49922
rect 53058 49870 53060 49922
rect 53004 49868 53060 49870
rect 53340 50370 53396 50372
rect 53340 50318 53342 50370
rect 53342 50318 53394 50370
rect 53394 50318 53396 50370
rect 53340 50316 53396 50318
rect 53452 50204 53508 50260
rect 53452 50034 53508 50036
rect 53452 49982 53454 50034
rect 53454 49982 53506 50034
rect 53506 49982 53508 50034
rect 53452 49980 53508 49982
rect 53116 49644 53172 49700
rect 53452 49644 53508 49700
rect 52892 48412 52948 48468
rect 53340 48748 53396 48804
rect 52780 47516 52836 47572
rect 53564 49250 53620 49252
rect 53564 49198 53566 49250
rect 53566 49198 53618 49250
rect 53618 49198 53620 49250
rect 53564 49196 53620 49198
rect 53788 48972 53844 49028
rect 53900 49756 53956 49812
rect 53676 48914 53732 48916
rect 53676 48862 53678 48914
rect 53678 48862 53730 48914
rect 53730 48862 53732 48914
rect 53676 48860 53732 48862
rect 53564 48802 53620 48804
rect 53564 48750 53566 48802
rect 53566 48750 53618 48802
rect 53618 48750 53620 48802
rect 53564 48748 53620 48750
rect 53900 48748 53956 48804
rect 54012 50316 54068 50372
rect 54012 48972 54068 49028
rect 53452 48524 53508 48580
rect 53788 48412 53844 48468
rect 53564 48076 53620 48132
rect 54124 48524 54180 48580
rect 54572 49026 54628 49028
rect 54572 48974 54574 49026
rect 54574 48974 54626 49026
rect 54626 48974 54628 49026
rect 54572 48972 54628 48974
rect 54236 48412 54292 48468
rect 54460 48860 54516 48916
rect 55132 50428 55188 50484
rect 55356 49698 55412 49700
rect 55356 49646 55358 49698
rect 55358 49646 55410 49698
rect 55410 49646 55412 49698
rect 55356 49644 55412 49646
rect 54796 48860 54852 48916
rect 55244 48860 55300 48916
rect 55356 48354 55412 48356
rect 55356 48302 55358 48354
rect 55358 48302 55410 48354
rect 55410 48302 55412 48354
rect 55356 48300 55412 48302
rect 53564 47292 53620 47348
rect 52220 46674 52276 46676
rect 52220 46622 52222 46674
rect 52222 46622 52274 46674
rect 52274 46622 52276 46674
rect 52220 46620 52276 46622
rect 51884 45500 51940 45556
rect 52108 45612 52164 45668
rect 52332 45890 52388 45892
rect 52332 45838 52334 45890
rect 52334 45838 52386 45890
rect 52386 45838 52388 45890
rect 52332 45836 52388 45838
rect 52668 46732 52724 46788
rect 52444 45500 52500 45556
rect 52668 45836 52724 45892
rect 52444 44492 52500 44548
rect 52220 44210 52276 44212
rect 52220 44158 52222 44210
rect 52222 44158 52274 44210
rect 52274 44158 52276 44210
rect 52220 44156 52276 44158
rect 52220 43708 52276 43764
rect 53116 46786 53172 46788
rect 53116 46734 53118 46786
rect 53118 46734 53170 46786
rect 53170 46734 53172 46786
rect 53116 46732 53172 46734
rect 53676 46898 53732 46900
rect 53676 46846 53678 46898
rect 53678 46846 53730 46898
rect 53730 46846 53732 46898
rect 53676 46844 53732 46846
rect 54460 47346 54516 47348
rect 54460 47294 54462 47346
rect 54462 47294 54514 47346
rect 54514 47294 54516 47346
rect 54460 47292 54516 47294
rect 55132 47628 55188 47684
rect 55132 47292 55188 47348
rect 55356 46844 55412 46900
rect 58044 57372 58100 57428
rect 58380 55356 58436 55412
rect 59724 57372 59780 57428
rect 59052 55132 59108 55188
rect 57932 53564 57988 53620
rect 58044 53228 58100 53284
rect 58044 52556 58100 52612
rect 58044 51212 58100 51268
rect 56140 49084 56196 49140
rect 56140 48860 56196 48916
rect 54908 46450 54964 46452
rect 54908 46398 54910 46450
rect 54910 46398 54962 46450
rect 54962 46398 54964 46450
rect 54908 46396 54964 46398
rect 53676 45890 53732 45892
rect 53676 45838 53678 45890
rect 53678 45838 53730 45890
rect 53730 45838 53732 45890
rect 53676 45836 53732 45838
rect 53004 44492 53060 44548
rect 53564 44098 53620 44100
rect 53564 44046 53566 44098
rect 53566 44046 53618 44098
rect 53618 44046 53620 44098
rect 53564 44044 53620 44046
rect 51660 43596 51716 43652
rect 51212 42082 51268 42084
rect 51212 42030 51214 42082
rect 51214 42030 51266 42082
rect 51266 42030 51268 42082
rect 51212 42028 51268 42030
rect 52556 43650 52612 43652
rect 52556 43598 52558 43650
rect 52558 43598 52610 43650
rect 52610 43598 52612 43650
rect 52556 43596 52612 43598
rect 53116 43708 53172 43764
rect 53564 43650 53620 43652
rect 53564 43598 53566 43650
rect 53566 43598 53618 43650
rect 53618 43598 53620 43650
rect 53564 43596 53620 43598
rect 51324 41916 51380 41972
rect 51660 41916 51716 41972
rect 52108 42028 52164 42084
rect 51100 41244 51156 41300
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50988 40796 51044 40852
rect 51324 41020 51380 41076
rect 50764 40740 50820 40742
rect 48636 40626 48692 40628
rect 48636 40574 48638 40626
rect 48638 40574 48690 40626
rect 48690 40574 48692 40626
rect 48636 40572 48692 40574
rect 49644 40572 49700 40628
rect 50764 40626 50820 40628
rect 50764 40574 50766 40626
rect 50766 40574 50818 40626
rect 50818 40574 50820 40626
rect 50764 40572 50820 40574
rect 48076 40348 48132 40404
rect 48412 40348 48468 40404
rect 49756 40348 49812 40404
rect 50316 40402 50372 40404
rect 50316 40350 50318 40402
rect 50318 40350 50370 40402
rect 50370 40350 50372 40402
rect 50316 40348 50372 40350
rect 50316 39730 50372 39732
rect 50316 39678 50318 39730
rect 50318 39678 50370 39730
rect 50370 39678 50372 39730
rect 50316 39676 50372 39678
rect 52332 41804 52388 41860
rect 53452 42588 53508 42644
rect 52780 42028 52836 42084
rect 52668 41410 52724 41412
rect 52668 41358 52670 41410
rect 52670 41358 52722 41410
rect 52722 41358 52724 41410
rect 52668 41356 52724 41358
rect 51548 40572 51604 40628
rect 51660 40796 51716 40852
rect 52220 40626 52276 40628
rect 52220 40574 52222 40626
rect 52222 40574 52274 40626
rect 52274 40574 52276 40626
rect 52220 40572 52276 40574
rect 52332 40348 52388 40404
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 44828 37436 44884 37492
rect 48300 37212 48356 37268
rect 53676 42642 53732 42644
rect 53676 42590 53678 42642
rect 53678 42590 53730 42642
rect 53730 42590 53732 42642
rect 53676 42588 53732 42590
rect 54460 44156 54516 44212
rect 54684 42812 54740 42868
rect 54236 42642 54292 42644
rect 54236 42590 54238 42642
rect 54238 42590 54290 42642
rect 54290 42590 54292 42642
rect 54236 42588 54292 42590
rect 54348 42476 54404 42532
rect 53676 41970 53732 41972
rect 53676 41918 53678 41970
rect 53678 41918 53730 41970
rect 53730 41918 53732 41970
rect 53676 41916 53732 41918
rect 53900 41858 53956 41860
rect 53900 41806 53902 41858
rect 53902 41806 53954 41858
rect 53954 41806 53956 41858
rect 53900 41804 53956 41806
rect 54124 41858 54180 41860
rect 54124 41806 54126 41858
rect 54126 41806 54178 41858
rect 54178 41806 54180 41858
rect 54124 41804 54180 41806
rect 53564 41692 53620 41748
rect 54572 41356 54628 41412
rect 55244 42476 55300 42532
rect 54796 41746 54852 41748
rect 54796 41694 54798 41746
rect 54798 41694 54850 41746
rect 54850 41694 54852 41746
rect 54796 41692 54852 41694
rect 52780 39676 52836 39732
rect 53452 40348 53508 40404
rect 52892 38722 52948 38724
rect 52892 38670 52894 38722
rect 52894 38670 52946 38722
rect 52946 38670 52948 38722
rect 52892 38668 52948 38670
rect 53676 38834 53732 38836
rect 53676 38782 53678 38834
rect 53678 38782 53730 38834
rect 53730 38782 53732 38834
rect 53676 38780 53732 38782
rect 54572 38780 54628 38836
rect 54236 38722 54292 38724
rect 54236 38670 54238 38722
rect 54238 38670 54290 38722
rect 54290 38670 54292 38722
rect 54236 38668 54292 38670
rect 57372 48466 57428 48468
rect 57372 48414 57374 48466
rect 57374 48414 57426 48466
rect 57426 48414 57428 48466
rect 57372 48412 57428 48414
rect 56252 47628 56308 47684
rect 56364 47516 56420 47572
rect 57260 47570 57316 47572
rect 57260 47518 57262 47570
rect 57262 47518 57314 47570
rect 57314 47518 57316 47570
rect 57260 47516 57316 47518
rect 58044 49138 58100 49140
rect 58044 49086 58046 49138
rect 58046 49086 58098 49138
rect 58098 49086 58100 49138
rect 58044 49084 58100 49086
rect 58044 47852 58100 47908
rect 57260 46396 57316 46452
rect 57484 46898 57540 46900
rect 57484 46846 57486 46898
rect 57486 46846 57538 46898
rect 57538 46846 57540 46898
rect 57484 46844 57540 46846
rect 58044 46508 58100 46564
rect 56364 45106 56420 45108
rect 56364 45054 56366 45106
rect 56366 45054 56418 45106
rect 56418 45054 56420 45106
rect 56364 45052 56420 45054
rect 56252 43596 56308 43652
rect 56252 42924 56308 42980
rect 56140 42812 56196 42868
rect 56364 42866 56420 42868
rect 56364 42814 56366 42866
rect 56366 42814 56418 42866
rect 56418 42814 56420 42866
rect 56364 42812 56420 42814
rect 55804 42476 55860 42532
rect 56812 42530 56868 42532
rect 56812 42478 56814 42530
rect 56814 42478 56866 42530
rect 56866 42478 56868 42530
rect 56812 42476 56868 42478
rect 56028 40908 56084 40964
rect 55244 38780 55300 38836
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 53564 37490 53620 37492
rect 53564 37438 53566 37490
rect 53566 37438 53618 37490
rect 53618 37438 53620 37490
rect 53564 37436 53620 37438
rect 54012 37436 54068 37492
rect 49532 37212 49588 37268
rect 42028 26290 42084 26292
rect 42028 26238 42030 26290
rect 42030 26238 42082 26290
rect 42082 26238 42084 26290
rect 42028 26236 42084 26238
rect 42812 26236 42868 26292
rect 47516 36482 47572 36484
rect 47516 36430 47518 36482
rect 47518 36430 47570 36482
rect 47570 36430 47572 36482
rect 47516 36428 47572 36430
rect 43932 25618 43988 25620
rect 43932 25566 43934 25618
rect 43934 25566 43986 25618
rect 43986 25566 43988 25618
rect 43932 25564 43988 25566
rect 43372 25228 43428 25284
rect 47516 25564 47572 25620
rect 43932 25228 43988 25284
rect 50876 36482 50932 36484
rect 50876 36430 50878 36482
rect 50878 36430 50930 36482
rect 50930 36430 50932 36482
rect 50876 36428 50932 36430
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 54348 35756 54404 35812
rect 54572 36428 54628 36484
rect 54572 35308 54628 35364
rect 54796 38668 54852 38724
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 56252 37100 56308 37156
rect 54908 36428 54964 36484
rect 56364 36428 56420 36484
rect 55244 36258 55300 36260
rect 55244 36206 55246 36258
rect 55246 36206 55298 36258
rect 55298 36206 55300 36258
rect 55244 36204 55300 36206
rect 55132 35308 55188 35364
rect 55132 23100 55188 23156
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 55804 36258 55860 36260
rect 55804 36206 55806 36258
rect 55806 36206 55858 36258
rect 55858 36206 55860 36258
rect 55804 36204 55860 36206
rect 55916 35756 55972 35812
rect 55356 35084 55412 35140
rect 56140 34972 56196 35028
rect 58044 45666 58100 45668
rect 58044 45614 58046 45666
rect 58046 45614 58098 45666
rect 58098 45614 58100 45666
rect 58044 45612 58100 45614
rect 57484 45052 57540 45108
rect 58044 44492 58100 44548
rect 57596 43650 57652 43652
rect 57596 43598 57598 43650
rect 57598 43598 57650 43650
rect 57650 43598 57652 43650
rect 57596 43596 57652 43598
rect 57932 43596 57988 43652
rect 57932 42812 57988 42868
rect 58044 40514 58100 40516
rect 58044 40462 58046 40514
rect 58046 40462 58098 40514
rect 58098 40462 58100 40514
rect 58044 40460 58100 40462
rect 58044 39116 58100 39172
rect 57372 37154 57428 37156
rect 57372 37102 57374 37154
rect 57374 37102 57426 37154
rect 57426 37102 57428 37154
rect 57372 37100 57428 37102
rect 58044 35026 58100 35028
rect 58044 34974 58046 35026
rect 58046 34974 58098 35026
rect 58098 34974 58100 35026
rect 58044 34972 58100 34974
rect 58044 31554 58100 31556
rect 58044 31502 58046 31554
rect 58046 31502 58098 31554
rect 58098 31502 58100 31554
rect 58044 31500 58100 31502
rect 57372 31052 57428 31108
rect 58044 30380 58100 30436
rect 58044 28418 58100 28420
rect 58044 28366 58046 28418
rect 58046 28366 58098 28418
rect 58098 28366 58100 28418
rect 58044 28364 58100 28366
rect 58044 24332 58100 24388
rect 57148 23100 57204 23156
rect 56252 22988 56308 23044
rect 57372 23042 57428 23044
rect 57372 22990 57374 23042
rect 57374 22990 57426 23042
rect 57426 22990 57428 23042
rect 57372 22988 57428 22990
rect 56252 19628 56308 19684
rect 57372 19628 57428 19684
rect 58044 15596 58100 15652
rect 58044 13580 58100 13636
rect 58044 10892 58100 10948
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 40908 3612 40964 3668
rect 58044 5516 58100 5572
rect 56252 4172 56308 4228
rect 57372 4226 57428 4228
rect 57372 4174 57374 4226
rect 57374 4174 57426 4226
rect 57426 4174 57428 4226
rect 57372 4172 57428 4174
rect 58044 3500 58100 3556
rect 28588 3442 28644 3444
rect 28588 3390 28590 3442
rect 28590 3390 28642 3442
rect 28642 3390 28644 3442
rect 28588 3388 28644 3390
rect 12908 3276 12964 3332
rect 13580 3330 13636 3332
rect 13580 3278 13582 3330
rect 13582 3278 13634 3330
rect 13634 3278 13636 3330
rect 13580 3276 13636 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 29372 3442 29428 3444
rect 29372 3390 29374 3442
rect 29374 3390 29426 3442
rect 29426 3390 29428 3442
rect 29372 3388 29428 3390
rect 36428 3276 36484 3332
rect 37100 3330 37156 3332
rect 37100 3278 37102 3330
rect 37102 3278 37154 3330
rect 37154 3278 37156 3330
rect 37100 3276 37156 3278
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 55916 2156 55972 2212
rect 58156 140 58212 196
<< metal3 >>
rect 200 59752 800 59976
rect 200 59080 800 59304
rect 59200 59080 59800 59304
rect 200 58436 800 58632
rect 59200 58436 59800 58632
rect 200 58408 3164 58436
rect 728 58380 3164 58408
rect 3220 58380 3230 58436
rect 57474 58380 57484 58436
rect 57540 58408 59800 58436
rect 57540 58380 59304 58408
rect 200 57736 800 57960
rect 59200 57736 59800 57960
rect 58034 57372 58044 57428
rect 58100 57372 59724 57428
rect 59780 57372 59790 57428
rect 200 57204 800 57288
rect 200 57148 4060 57204
rect 4116 57148 4126 57204
rect 200 57064 800 57148
rect 59200 57064 59800 57288
rect 200 56392 800 56616
rect 56578 56588 56588 56644
rect 56644 56588 57372 56644
rect 57428 56588 57438 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 59200 56392 59800 56616
rect 36418 56252 36428 56308
rect 36484 56252 37100 56308
rect 37156 56252 37166 56308
rect 46498 56252 46508 56308
rect 46564 56252 47964 56308
rect 48020 56252 48030 56308
rect 12786 56028 12796 56084
rect 12852 56028 15036 56084
rect 15092 56028 15102 56084
rect 200 55720 800 55944
rect 46274 55916 46284 55972
rect 46340 55916 47180 55972
rect 47236 55916 47246 55972
rect 55906 55916 55916 55972
rect 55972 55916 57260 55972
rect 57316 55916 57326 55972
rect 59200 55720 59800 55944
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 54002 55356 54012 55412
rect 54068 55356 55020 55412
rect 55076 55356 58380 55412
rect 58436 55356 58446 55412
rect 728 55272 1820 55300
rect 200 55244 1820 55272
rect 1876 55244 1886 55300
rect 3042 55244 3052 55300
rect 3108 55244 3724 55300
rect 3780 55244 3790 55300
rect 200 55048 800 55244
rect 12898 55132 12908 55188
rect 12964 55132 13692 55188
rect 13748 55132 13758 55188
rect 56242 55132 56252 55188
rect 56308 55132 56700 55188
rect 56756 55132 59052 55188
rect 59108 55132 59118 55188
rect 59200 55048 59800 55272
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 1474 54684 1484 54740
rect 1540 54684 2492 54740
rect 2548 54684 2558 54740
rect 48850 54684 48860 54740
rect 48916 54684 50540 54740
rect 50596 54684 50606 54740
rect 728 54600 1932 54628
rect 200 54572 1932 54600
rect 1988 54572 1998 54628
rect 52210 54572 52220 54628
rect 52276 54572 53564 54628
rect 53620 54572 53630 54628
rect 200 54376 800 54572
rect 15026 54348 15036 54404
rect 15092 54348 41580 54404
rect 41636 54348 41646 54404
rect 44482 54348 44492 54404
rect 44548 54348 44940 54404
rect 44996 54348 45612 54404
rect 45668 54348 45678 54404
rect 59200 54376 59800 54600
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 728 53928 1820 53956
rect 200 53900 1820 53928
rect 1876 53900 1886 53956
rect 200 53704 800 53900
rect 45602 53788 45612 53844
rect 45668 53788 47292 53844
rect 47348 53788 47358 53844
rect 44706 53676 44716 53732
rect 44772 53676 51884 53732
rect 51940 53676 51950 53732
rect 59200 53704 59800 53928
rect 47282 53564 47292 53620
rect 47348 53564 50540 53620
rect 50596 53564 57932 53620
rect 57988 53564 57998 53620
rect 7186 53452 7196 53508
rect 7252 53452 46732 53508
rect 46788 53452 47964 53508
rect 48020 53452 48030 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 728 53256 1932 53284
rect 200 53228 1932 53256
rect 1988 53228 1998 53284
rect 58034 53228 58044 53284
rect 58100 53256 59304 53284
rect 58100 53228 59800 53256
rect 200 53032 800 53228
rect 44146 53116 44156 53172
rect 44212 53116 44380 53172
rect 44436 53116 45276 53172
rect 45332 53116 45342 53172
rect 44818 53004 44828 53060
rect 44884 53004 45500 53060
rect 45556 53004 45566 53060
rect 48066 53004 48076 53060
rect 48132 53004 49420 53060
rect 49476 53004 49486 53060
rect 59200 53032 59800 53228
rect 44706 52892 44716 52948
rect 44772 52892 45612 52948
rect 45668 52892 45678 52948
rect 3714 52780 3724 52836
rect 3780 52780 50092 52836
rect 50148 52780 50158 52836
rect 51650 52780 51660 52836
rect 51716 52780 52220 52836
rect 52276 52780 52286 52836
rect 728 52584 1820 52612
rect 200 52556 1820 52584
rect 1876 52556 1886 52612
rect 58034 52556 58044 52612
rect 58100 52584 59304 52612
rect 58100 52556 59800 52584
rect 200 52360 800 52556
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 59200 52360 59800 52556
rect 42802 52220 42812 52276
rect 42868 52220 43260 52276
rect 43316 52220 44492 52276
rect 44548 52220 44558 52276
rect 55122 52220 55132 52276
rect 55188 52220 55580 52276
rect 55636 52220 55646 52276
rect 3490 51996 3500 52052
rect 3556 51996 39900 52052
rect 39956 51996 39966 52052
rect 46722 51996 46732 52052
rect 46788 51996 47292 52052
rect 47348 51996 47358 52052
rect 44034 51884 44044 51940
rect 44100 51884 44716 51940
rect 44772 51884 44782 51940
rect 45714 51884 45724 51940
rect 45780 51884 46396 51940
rect 46452 51884 46462 51940
rect 48178 51884 48188 51940
rect 48244 51884 48748 51940
rect 48804 51884 48814 51940
rect 48962 51884 48972 51940
rect 49028 51884 49644 51940
rect 49700 51884 49710 51940
rect 45724 51828 45780 51884
rect 44818 51772 44828 51828
rect 44884 51772 45780 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 46386 51660 46396 51716
rect 46452 51660 48636 51716
rect 48692 51660 48972 51716
rect 49028 51660 49038 51716
rect 48290 51548 48300 51604
rect 48356 51548 49420 51604
rect 49476 51548 49486 51604
rect 44034 51436 44044 51492
rect 44100 51436 44828 51492
rect 44884 51436 44894 51492
rect 45826 51436 45836 51492
rect 45892 51436 48188 51492
rect 48244 51436 48254 51492
rect 49634 51436 49644 51492
rect 49700 51436 50652 51492
rect 50708 51436 50718 51492
rect 44594 51324 44604 51380
rect 44660 51324 45948 51380
rect 46004 51324 46396 51380
rect 46452 51324 46462 51380
rect 728 51240 1820 51268
rect 200 51212 1820 51240
rect 1876 51212 1886 51268
rect 49746 51212 49756 51268
rect 49812 51212 50204 51268
rect 50260 51212 50270 51268
rect 58034 51212 58044 51268
rect 58100 51240 59304 51268
rect 58100 51212 59800 51240
rect 200 51016 800 51212
rect 41682 50988 41692 51044
rect 41748 50988 48188 51044
rect 48244 50988 48254 51044
rect 59200 51016 59800 51212
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 4834 50652 4844 50708
rect 4900 50652 39564 50708
rect 39620 50652 39630 50708
rect 46274 50652 46284 50708
rect 46340 50652 46732 50708
rect 46788 50652 46798 50708
rect 200 50344 800 50568
rect 45378 50540 45388 50596
rect 45444 50540 48748 50596
rect 48804 50540 49308 50596
rect 49364 50540 49756 50596
rect 49812 50540 49822 50596
rect 44706 50428 44716 50484
rect 44772 50428 45276 50484
rect 45332 50428 45342 50484
rect 47282 50428 47292 50484
rect 47348 50428 47964 50484
rect 48020 50428 48636 50484
rect 48692 50428 48702 50484
rect 50642 50428 50652 50484
rect 50708 50428 52780 50484
rect 52836 50428 55132 50484
rect 55188 50428 55198 50484
rect 48514 50316 48524 50372
rect 48580 50316 50876 50372
rect 50932 50316 52108 50372
rect 52164 50316 53340 50372
rect 53396 50316 54012 50372
rect 54068 50316 54078 50372
rect 59200 50344 59800 50568
rect 52994 50204 53004 50260
rect 53060 50204 53452 50260
rect 53508 50204 53518 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 51874 50092 51884 50148
rect 51940 50092 52556 50148
rect 52612 50092 52622 50148
rect 46386 49980 46396 50036
rect 46452 49980 47404 50036
rect 47460 49980 47470 50036
rect 51762 49980 51772 50036
rect 51828 49980 53452 50036
rect 53508 49980 53518 50036
rect 200 49672 800 49896
rect 49634 49868 49644 49924
rect 49700 49868 53004 49924
rect 53060 49868 53070 49924
rect 44258 49756 44268 49812
rect 44324 49756 44604 49812
rect 44660 49756 44670 49812
rect 44930 49756 44940 49812
rect 44996 49756 45612 49812
rect 45668 49756 45678 49812
rect 47954 49756 47964 49812
rect 48020 49756 48412 49812
rect 48468 49756 48478 49812
rect 48626 49756 48636 49812
rect 48692 49756 49532 49812
rect 49588 49756 50988 49812
rect 51044 49756 51324 49812
rect 51380 49756 51772 49812
rect 51828 49756 53900 49812
rect 53956 49756 53966 49812
rect 59200 49700 59800 49896
rect 48850 49644 48860 49700
rect 48916 49644 48926 49700
rect 49970 49644 49980 49700
rect 50036 49644 51548 49700
rect 51604 49644 53116 49700
rect 53172 49644 53452 49700
rect 53508 49644 53518 49700
rect 55346 49644 55356 49700
rect 55412 49672 59800 49700
rect 55412 49644 59304 49672
rect 48860 49588 48916 49644
rect 48860 49532 49084 49588
rect 49140 49532 49150 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 50306 49308 50316 49364
rect 50372 49308 51996 49364
rect 52052 49308 52062 49364
rect 200 49000 800 49224
rect 52658 49196 52668 49252
rect 52724 49196 53564 49252
rect 53620 49196 53630 49252
rect 42690 49084 42700 49140
rect 42756 49084 44268 49140
rect 44324 49084 44334 49140
rect 48738 49084 48748 49140
rect 48804 49084 50092 49140
rect 50148 49084 50158 49140
rect 56130 49084 56140 49140
rect 56196 49084 58044 49140
rect 58100 49084 58110 49140
rect 44482 48972 44492 49028
rect 44548 48972 45500 49028
rect 45556 48972 45566 49028
rect 45826 48972 45836 49028
rect 45892 48972 46508 49028
rect 46564 48972 47180 49028
rect 47236 48972 47246 49028
rect 48514 48972 48524 49028
rect 48580 48972 49868 49028
rect 49924 48972 49934 49028
rect 51650 48972 51660 49028
rect 51716 48972 52220 49028
rect 52276 48972 52286 49028
rect 52546 48972 52556 49028
rect 52612 48972 53788 49028
rect 53844 48972 53854 49028
rect 54002 48972 54012 49028
rect 54068 48972 54572 49028
rect 54628 48972 54638 49028
rect 59200 49000 59800 49224
rect 44146 48860 44156 48916
rect 44212 48860 45948 48916
rect 46004 48860 46014 48916
rect 46946 48860 46956 48916
rect 47012 48860 47404 48916
rect 47460 48860 49756 48916
rect 49812 48860 49822 48916
rect 50194 48860 50204 48916
rect 50260 48860 50540 48916
rect 50596 48860 50876 48916
rect 50932 48860 50942 48916
rect 51548 48860 53676 48916
rect 53732 48860 54460 48916
rect 54516 48860 54526 48916
rect 54786 48860 54796 48916
rect 54852 48860 55244 48916
rect 55300 48860 56140 48916
rect 56196 48860 56206 48916
rect 47170 48748 47180 48804
rect 47236 48748 47516 48804
rect 47572 48748 49196 48804
rect 49252 48748 49262 48804
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 51548 48580 51604 48860
rect 53330 48748 53340 48804
rect 53396 48748 53564 48804
rect 53620 48748 53900 48804
rect 53956 48748 53966 48804
rect 52742 48636 52780 48692
rect 52836 48636 52846 48692
rect 200 48328 800 48552
rect 46386 48524 46396 48580
rect 46452 48524 47628 48580
rect 47684 48524 47694 48580
rect 51538 48524 51548 48580
rect 51604 48524 51614 48580
rect 53442 48524 53452 48580
rect 53508 48524 54124 48580
rect 54180 48524 54190 48580
rect 49858 48412 49868 48468
rect 49924 48412 52108 48468
rect 52164 48412 52892 48468
rect 52948 48412 53788 48468
rect 53844 48412 54236 48468
rect 54292 48412 57372 48468
rect 57428 48412 57438 48468
rect 59200 48356 59800 48552
rect 47058 48300 47068 48356
rect 47124 48300 47516 48356
rect 47572 48300 48300 48356
rect 48356 48300 48366 48356
rect 55346 48300 55356 48356
rect 55412 48328 59800 48356
rect 55412 48300 59304 48328
rect 46386 48188 46396 48244
rect 46452 48188 46732 48244
rect 46788 48188 47292 48244
rect 47348 48188 47358 48244
rect 50418 48076 50428 48132
rect 50484 48076 50988 48132
rect 51044 48076 53564 48132
rect 53620 48076 53630 48132
rect 200 47656 800 47880
rect 58034 47852 58044 47908
rect 58100 47880 59304 47908
rect 58100 47852 59800 47880
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 43250 47628 43260 47684
rect 43316 47628 44268 47684
rect 44324 47628 44334 47684
rect 55122 47628 55132 47684
rect 55188 47628 56252 47684
rect 56308 47628 56318 47684
rect 59200 47656 59800 47852
rect 43138 47516 43148 47572
rect 43204 47516 44380 47572
rect 44436 47516 45500 47572
rect 45556 47516 45566 47572
rect 49746 47516 49756 47572
rect 49812 47516 49980 47572
rect 50036 47516 50652 47572
rect 50708 47516 51212 47572
rect 51268 47516 52780 47572
rect 52836 47516 52846 47572
rect 56354 47516 56364 47572
rect 56420 47516 57260 47572
rect 57316 47516 57326 47572
rect 46162 47404 46172 47460
rect 46228 47404 47068 47460
rect 47124 47404 47134 47460
rect 53554 47292 53564 47348
rect 53620 47292 54460 47348
rect 54516 47292 55132 47348
rect 55188 47292 55198 47348
rect 728 47208 1820 47236
rect 200 47180 1820 47208
rect 1876 47180 1886 47236
rect 43362 47180 43372 47236
rect 43428 47180 44268 47236
rect 44324 47180 46396 47236
rect 46452 47180 46462 47236
rect 200 46984 800 47180
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 48290 46956 48300 47012
rect 48356 46956 48748 47012
rect 48804 46956 49308 47012
rect 49364 46956 49532 47012
rect 49588 46956 50204 47012
rect 50260 46956 50270 47012
rect 50978 46956 50988 47012
rect 51044 46956 51436 47012
rect 51492 46956 51502 47012
rect 59200 46984 59800 47208
rect 48178 46844 48188 46900
rect 48244 46844 49980 46900
rect 50036 46844 50046 46900
rect 51090 46844 51100 46900
rect 51156 46844 51548 46900
rect 51604 46844 53676 46900
rect 53732 46844 53742 46900
rect 55346 46844 55356 46900
rect 55412 46844 57484 46900
rect 57540 46844 57550 46900
rect 46162 46732 46172 46788
rect 46228 46732 46732 46788
rect 46788 46732 47068 46788
rect 47124 46732 47134 46788
rect 52658 46732 52668 46788
rect 52724 46732 53116 46788
rect 53172 46732 53182 46788
rect 43026 46620 43036 46676
rect 43092 46620 46508 46676
rect 46564 46620 46956 46676
rect 47012 46620 47292 46676
rect 47348 46620 48524 46676
rect 48580 46620 48860 46676
rect 48916 46620 48926 46676
rect 51986 46620 51996 46676
rect 52052 46620 52220 46676
rect 52276 46620 52286 46676
rect 200 46312 800 46536
rect 58034 46508 58044 46564
rect 58100 46536 59304 46564
rect 58100 46508 59800 46536
rect 47506 46396 47516 46452
rect 47572 46396 49644 46452
rect 49700 46396 51884 46452
rect 51940 46396 51950 46452
rect 54898 46396 54908 46452
rect 54964 46396 57260 46452
rect 57316 46396 57326 46452
rect 47058 46284 47068 46340
rect 47124 46284 47628 46340
rect 47684 46284 47694 46340
rect 59200 46312 59800 46508
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 48738 45948 48748 46004
rect 48804 45948 50092 46004
rect 50148 45948 50764 46004
rect 50820 45948 50830 46004
rect 200 45668 800 45864
rect 48178 45836 48188 45892
rect 48244 45836 49644 45892
rect 49700 45836 49710 45892
rect 51314 45836 51324 45892
rect 51380 45836 52332 45892
rect 52388 45836 52398 45892
rect 52658 45836 52668 45892
rect 52724 45836 53676 45892
rect 53732 45836 53742 45892
rect 42690 45724 42700 45780
rect 42756 45724 43148 45780
rect 43204 45724 47068 45780
rect 47124 45724 47134 45780
rect 48402 45724 48412 45780
rect 48468 45724 49196 45780
rect 49252 45724 49262 45780
rect 59200 45668 59800 45864
rect 200 45640 2492 45668
rect 728 45612 2492 45640
rect 2548 45612 2558 45668
rect 48626 45612 48636 45668
rect 48692 45612 49644 45668
rect 49700 45612 50988 45668
rect 51044 45612 51054 45668
rect 51314 45612 51324 45668
rect 51380 45612 52108 45668
rect 52164 45612 52174 45668
rect 58034 45612 58044 45668
rect 58100 45640 59800 45668
rect 58100 45612 59304 45640
rect 50988 45556 51044 45612
rect 50988 45500 51436 45556
rect 51492 45500 51502 45556
rect 51874 45500 51884 45556
rect 51940 45500 52444 45556
rect 52500 45500 52510 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 46722 45388 46732 45444
rect 46788 45388 48972 45444
rect 49028 45388 49038 45444
rect 728 45192 1708 45220
rect 200 45164 1708 45192
rect 1764 45164 1774 45220
rect 42802 45164 42812 45220
rect 42868 45164 43596 45220
rect 43652 45164 43662 45220
rect 200 44968 800 45164
rect 44258 45052 44268 45108
rect 44324 45052 45052 45108
rect 45108 45052 45118 45108
rect 46498 45052 46508 45108
rect 46564 45052 48188 45108
rect 48244 45052 48254 45108
rect 56354 45052 56364 45108
rect 56420 45052 57484 45108
rect 57540 45052 57550 45108
rect 44482 44940 44492 44996
rect 44548 44940 46060 44996
rect 46116 44940 47964 44996
rect 48020 44940 48030 44996
rect 59200 44968 59800 45192
rect 44706 44828 44716 44884
rect 44772 44828 45836 44884
rect 45892 44828 48524 44884
rect 48580 44828 48590 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 728 44520 1820 44548
rect 200 44492 1820 44520
rect 1876 44492 1886 44548
rect 52434 44492 52444 44548
rect 52500 44492 53004 44548
rect 53060 44492 53070 44548
rect 58034 44492 58044 44548
rect 58100 44520 59304 44548
rect 58100 44492 59800 44520
rect 200 44296 800 44492
rect 43698 44380 43708 44436
rect 43764 44380 45500 44436
rect 45556 44380 45566 44436
rect 44594 44268 44604 44324
rect 44660 44268 45948 44324
rect 46004 44268 46014 44324
rect 59200 44296 59800 44492
rect 43474 44156 43484 44212
rect 43540 44156 44100 44212
rect 48738 44156 48748 44212
rect 48804 44156 52220 44212
rect 52276 44156 54460 44212
rect 54516 44156 54526 44212
rect 44044 44100 44100 44156
rect 44034 44044 44044 44100
rect 44100 44044 45052 44100
rect 45108 44044 53564 44100
rect 53620 44044 53630 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 200 43624 800 43848
rect 52210 43708 52220 43764
rect 52276 43708 53116 43764
rect 53172 43708 53182 43764
rect 51202 43596 51212 43652
rect 51268 43596 51660 43652
rect 51716 43596 52556 43652
rect 52612 43596 53564 43652
rect 53620 43596 53630 43652
rect 56242 43596 56252 43652
rect 56308 43596 57596 43652
rect 57652 43596 57932 43652
rect 57988 43596 57998 43652
rect 59200 43624 59800 43848
rect 48962 43372 48972 43428
rect 49028 43372 50876 43428
rect 50932 43372 51100 43428
rect 51156 43372 51166 43428
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 43652 42924 44940 42980
rect 44996 42924 56252 42980
rect 56308 42924 56318 42980
rect 40114 42700 40124 42756
rect 40180 42700 42028 42756
rect 42084 42700 43596 42756
rect 43652 42700 43708 42924
rect 45378 42812 45388 42868
rect 45444 42812 46284 42868
rect 46340 42812 46350 42868
rect 48514 42812 48524 42868
rect 48580 42812 49420 42868
rect 49476 42812 49868 42868
rect 49924 42812 49934 42868
rect 54674 42812 54684 42868
rect 54740 42812 56140 42868
rect 56196 42812 56364 42868
rect 56420 42812 57932 42868
rect 57988 42812 57998 42868
rect 39442 42588 39452 42644
rect 39508 42588 40796 42644
rect 40852 42588 40862 42644
rect 53442 42588 53452 42644
rect 53508 42588 53676 42644
rect 53732 42588 54236 42644
rect 54292 42588 54302 42644
rect 200 42280 800 42504
rect 46162 42476 46172 42532
rect 46228 42476 46732 42532
rect 46788 42476 46798 42532
rect 48290 42476 48300 42532
rect 48356 42476 50988 42532
rect 51044 42476 54348 42532
rect 54404 42476 54414 42532
rect 55234 42476 55244 42532
rect 55300 42476 55804 42532
rect 55860 42476 56812 42532
rect 56868 42476 56878 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 59200 42280 59800 42504
rect 51202 42028 51212 42084
rect 51268 42028 52108 42084
rect 52164 42028 52174 42084
rect 52770 42028 52780 42084
rect 52836 42028 54180 42084
rect 46386 41916 46396 41972
rect 46452 41916 48076 41972
rect 48132 41916 48142 41972
rect 49746 41916 49756 41972
rect 49812 41916 50428 41972
rect 50484 41916 51324 41972
rect 51380 41916 51390 41972
rect 51650 41916 51660 41972
rect 51716 41916 53676 41972
rect 53732 41916 53742 41972
rect 54124 41860 54180 42028
rect 200 41608 800 41832
rect 48626 41804 48636 41860
rect 48692 41804 49532 41860
rect 49588 41804 49598 41860
rect 52322 41804 52332 41860
rect 52388 41804 53900 41860
rect 53956 41804 53966 41860
rect 54114 41804 54124 41860
rect 54180 41804 54190 41860
rect 47954 41692 47964 41748
rect 48020 41692 49980 41748
rect 50036 41692 50316 41748
rect 50372 41692 50876 41748
rect 50932 41692 50942 41748
rect 53554 41692 53564 41748
rect 53620 41692 54796 41748
rect 54852 41692 54862 41748
rect 59200 41608 59800 41832
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 46610 41356 46620 41412
rect 46676 41356 47404 41412
rect 47460 41356 47470 41412
rect 48066 41356 48076 41412
rect 48132 41356 49644 41412
rect 49700 41356 49710 41412
rect 52658 41356 52668 41412
rect 52724 41356 54572 41412
rect 54628 41356 54638 41412
rect 48402 41244 48412 41300
rect 48468 41244 51100 41300
rect 51156 41244 51166 41300
rect 200 40964 800 41160
rect 46610 41132 46620 41188
rect 46676 41132 46844 41188
rect 46900 41132 47292 41188
rect 47348 41132 47358 41188
rect 48290 41132 48300 41188
rect 48356 41132 49700 41188
rect 49644 41076 49700 41132
rect 46386 41020 46396 41076
rect 46452 41020 47404 41076
rect 47460 41020 48188 41076
rect 48244 41020 48254 41076
rect 49634 41020 49644 41076
rect 49700 41020 50204 41076
rect 50260 41020 51324 41076
rect 51380 41020 51390 41076
rect 59200 40964 59800 41160
rect 200 40936 2492 40964
rect 728 40908 2492 40936
rect 2548 40908 2558 40964
rect 56018 40908 56028 40964
rect 56084 40936 59800 40964
rect 56084 40908 59304 40936
rect 50978 40796 50988 40852
rect 51044 40796 51660 40852
rect 51716 40796 51726 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 44482 40572 44492 40628
rect 44548 40572 45276 40628
rect 45332 40572 46284 40628
rect 46340 40572 47068 40628
rect 47124 40572 47964 40628
rect 48020 40572 48636 40628
rect 48692 40572 48702 40628
rect 49634 40572 49644 40628
rect 49700 40572 50764 40628
rect 50820 40572 50830 40628
rect 51538 40572 51548 40628
rect 51604 40572 52220 40628
rect 52276 40572 52286 40628
rect 728 40488 1708 40516
rect 200 40460 1708 40488
rect 1764 40460 1774 40516
rect 46946 40460 46956 40516
rect 47012 40460 47404 40516
rect 47460 40460 47852 40516
rect 47908 40460 47918 40516
rect 58034 40460 58044 40516
rect 58100 40488 59304 40516
rect 58100 40460 59800 40488
rect 200 40264 800 40460
rect 40898 40348 40908 40404
rect 40964 40348 42364 40404
rect 42420 40348 42430 40404
rect 48066 40348 48076 40404
rect 48132 40348 48412 40404
rect 48468 40348 49756 40404
rect 49812 40348 50316 40404
rect 50372 40348 52332 40404
rect 52388 40348 53452 40404
rect 53508 40348 53518 40404
rect 59200 40264 59800 40460
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 728 39816 1820 39844
rect 200 39788 1820 39816
rect 1876 39788 1886 39844
rect 200 39592 800 39788
rect 50306 39676 50316 39732
rect 50372 39676 52780 39732
rect 52836 39676 52846 39732
rect 59200 39592 59800 39816
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 728 39144 1820 39172
rect 200 39116 1820 39144
rect 1876 39116 1886 39172
rect 58034 39116 58044 39172
rect 58100 39144 59304 39172
rect 58100 39116 59800 39144
rect 200 38920 800 39116
rect 59200 38920 59800 39116
rect 53666 38780 53676 38836
rect 53732 38780 54572 38836
rect 54628 38780 55244 38836
rect 55300 38780 55310 38836
rect 52882 38668 52892 38724
rect 52948 38668 54236 38724
rect 54292 38668 54796 38724
rect 54852 38668 54862 38724
rect 200 38248 800 38472
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 59200 38248 59800 38472
rect 200 37576 800 37800
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 59200 37576 59800 37800
rect 44818 37436 44828 37492
rect 44884 37436 53564 37492
rect 53620 37436 54012 37492
rect 54068 37436 54078 37492
rect 48290 37212 48300 37268
rect 48356 37212 49532 37268
rect 49588 37212 49598 37268
rect 200 36904 800 37128
rect 56242 37100 56252 37156
rect 56308 37100 57372 37156
rect 57428 37128 59304 37156
rect 57428 37100 59800 37128
rect 59200 36904 59800 37100
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 200 36232 800 36456
rect 47506 36428 47516 36484
rect 47572 36428 50876 36484
rect 50932 36428 54572 36484
rect 54628 36428 54908 36484
rect 54964 36428 56364 36484
rect 56420 36428 56430 36484
rect 55234 36204 55244 36260
rect 55300 36204 55804 36260
rect 55860 36204 55870 36260
rect 59200 36232 59800 36456
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 200 35560 800 35784
rect 54338 35756 54348 35812
rect 54404 35756 55916 35812
rect 55972 35756 55982 35812
rect 59200 35560 59800 35784
rect 54562 35308 54572 35364
rect 54628 35308 55132 35364
rect 55188 35308 55198 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 728 35112 1820 35140
rect 200 35084 1820 35112
rect 1876 35084 1886 35140
rect 55346 35084 55356 35140
rect 55412 35112 59304 35140
rect 55412 35084 59800 35112
rect 200 34888 800 35084
rect 56130 34972 56140 35028
rect 56196 34972 58044 35028
rect 58100 34972 58110 35028
rect 59200 34888 59800 35084
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 200 33544 800 33768
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 59200 33544 59800 33768
rect 200 32872 800 33096
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 59200 32872 59800 33096
rect 200 32200 800 32424
rect 59200 32200 59800 32424
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 200 31556 800 31752
rect 59200 31556 59800 31752
rect 200 31528 1820 31556
rect 728 31500 1820 31528
rect 1876 31500 1886 31556
rect 58034 31500 58044 31556
rect 58100 31528 59800 31556
rect 58100 31500 59304 31528
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 728 31080 2492 31108
rect 200 31052 2492 31080
rect 2548 31052 2558 31108
rect 57362 31052 57372 31108
rect 57428 31080 59304 31108
rect 57428 31052 59800 31080
rect 200 30856 800 31052
rect 59200 30856 59800 31052
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 200 30184 800 30408
rect 58034 30380 58044 30436
rect 58100 30408 59304 30436
rect 58100 30380 59800 30408
rect 59200 30184 59800 30380
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 200 29512 800 29736
rect 59200 29512 59800 29736
rect 200 28840 800 29064
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 59200 28840 59800 29064
rect 728 28392 1820 28420
rect 200 28364 1820 28392
rect 1876 28364 1886 28420
rect 58034 28364 58044 28420
rect 58100 28392 59304 28420
rect 58100 28364 59800 28392
rect 200 28168 800 28364
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 59200 28168 59800 28364
rect 200 27496 800 27720
rect 59200 27496 59800 27720
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 200 26964 800 27048
rect 200 26908 1820 26964
rect 1876 26908 1886 26964
rect 200 26824 800 26908
rect 59200 26824 59800 27048
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 200 26152 800 26376
rect 42018 26236 42028 26292
rect 42084 26236 42812 26292
rect 42868 26236 42878 26292
rect 59200 26152 59800 26376
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 43922 25564 43932 25620
rect 43988 25564 47516 25620
rect 47572 25564 47582 25620
rect 3042 25228 3052 25284
rect 3108 25228 3612 25284
rect 3668 25228 40460 25284
rect 40516 25228 40526 25284
rect 43362 25228 43372 25284
rect 43428 25228 43932 25284
rect 43988 25228 43998 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 728 25032 1932 25060
rect 200 25004 1932 25032
rect 1988 25004 1998 25060
rect 200 24808 800 25004
rect 59200 24808 59800 25032
rect 200 24136 800 24360
rect 58034 24332 58044 24388
rect 58100 24360 59304 24388
rect 58100 24332 59800 24360
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 59200 24136 59800 24332
rect 200 23464 800 23688
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 59200 23464 59800 23688
rect 55122 23100 55132 23156
rect 55188 23100 57148 23156
rect 57204 23100 57214 23156
rect 728 23016 1820 23044
rect 200 22988 1820 23016
rect 1876 22988 1886 23044
rect 56242 22988 56252 23044
rect 56308 22988 57372 23044
rect 57428 23016 59304 23044
rect 57428 22988 59800 23016
rect 200 22792 800 22988
rect 59200 22792 59800 22988
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 200 22120 800 22344
rect 59200 22120 59800 22344
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 728 21672 1708 21700
rect 200 21644 1708 21672
rect 1764 21644 1774 21700
rect 200 21448 800 21644
rect 59200 21448 59800 21672
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 728 21000 1820 21028
rect 200 20972 1820 21000
rect 1876 20972 1886 21028
rect 200 20776 800 20972
rect 59200 20776 59800 21000
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 200 20104 800 20328
rect 59200 20104 59800 20328
rect 728 19656 1820 19684
rect 200 19628 1820 19656
rect 1876 19628 1886 19684
rect 56242 19628 56252 19684
rect 56308 19628 57372 19684
rect 57428 19656 59304 19684
rect 57428 19628 59800 19656
rect 200 19432 800 19628
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 59200 19432 59800 19628
rect 200 18760 800 18984
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 59200 18760 59800 18984
rect 728 18312 1820 18340
rect 200 18284 1820 18312
rect 1876 18284 1886 18340
rect 200 18088 800 18284
rect 59200 18088 59800 18312
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 200 17416 800 17640
rect 59200 17416 59800 17640
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 728 16296 1820 16324
rect 200 16268 1820 16296
rect 1876 16268 1886 16324
rect 200 16072 800 16268
rect 59200 16072 59800 16296
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 200 15400 800 15624
rect 58034 15596 58044 15652
rect 58100 15624 59304 15652
rect 58100 15596 59800 15624
rect 59200 15400 59800 15596
rect 728 14952 1820 14980
rect 200 14924 1820 14952
rect 1876 14924 1886 14980
rect 200 14728 800 14924
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 59200 14728 59800 14952
rect 728 14280 1820 14308
rect 200 14252 1820 14280
rect 1876 14252 1886 14308
rect 200 14056 800 14252
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 59200 14056 59800 14280
rect 200 13384 800 13608
rect 58034 13580 58044 13636
rect 58100 13608 59304 13636
rect 58100 13580 59800 13608
rect 59200 13384 59800 13580
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 200 12740 800 12936
rect 200 12712 1820 12740
rect 728 12684 1820 12712
rect 1876 12684 1886 12740
rect 59200 12712 59800 12936
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 200 12040 800 12264
rect 59200 12040 59800 12264
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 200 11368 800 11592
rect 59200 11368 59800 11592
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 200 10696 800 10920
rect 58034 10892 58044 10948
rect 58100 10920 59304 10948
rect 58100 10892 59800 10920
rect 59200 10696 59800 10892
rect 728 10248 1820 10276
rect 200 10220 1820 10248
rect 1876 10220 1886 10276
rect 200 10024 800 10220
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 59200 10024 59800 10248
rect 728 9576 1820 9604
rect 200 9548 1820 9576
rect 1876 9548 1886 9604
rect 200 9352 800 9548
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 59200 9352 59800 9576
rect 200 8680 800 8904
rect 59200 8680 59800 8904
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 200 7336 800 7560
rect 59200 7336 59800 7560
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 200 6664 800 6888
rect 59200 6664 59800 6888
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 728 6216 1820 6244
rect 200 6188 1820 6216
rect 1876 6188 1886 6244
rect 200 5992 800 6188
rect 59200 5992 59800 6216
rect 200 5320 800 5544
rect 58034 5516 58044 5572
rect 58100 5544 59304 5572
rect 58100 5516 59800 5544
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 59200 5320 59800 5516
rect 728 4872 1820 4900
rect 200 4844 1820 4872
rect 1876 4844 1886 4900
rect 200 4648 800 4844
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 59200 4648 59800 4872
rect 200 3976 800 4200
rect 11554 4172 11564 4228
rect 11620 4172 13020 4228
rect 13076 4172 13086 4228
rect 56242 4172 56252 4228
rect 56308 4172 57372 4228
rect 57428 4200 59304 4228
rect 57428 4172 59800 4200
rect 59200 3976 59800 4172
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 30706 3724 30716 3780
rect 30772 3724 39452 3780
rect 39508 3724 39518 3780
rect 12786 3612 12796 3668
rect 12852 3612 40908 3668
rect 40964 3612 40974 3668
rect 200 3304 800 3528
rect 58034 3500 58044 3556
rect 58100 3528 59304 3556
rect 58100 3500 59800 3528
rect 28578 3388 28588 3444
rect 28644 3388 29372 3444
rect 29428 3388 29438 3444
rect 12898 3276 12908 3332
rect 12964 3276 13580 3332
rect 13636 3276 13646 3332
rect 36418 3276 36428 3332
rect 36484 3276 37100 3332
rect 37156 3276 37166 3332
rect 59200 3304 59800 3500
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 200 2632 800 2856
rect 59200 2632 59800 2856
rect 728 2184 1932 2212
rect 200 2156 1932 2184
rect 1988 2156 1998 2212
rect 55906 2156 55916 2212
rect 55972 2184 59304 2212
rect 55972 2156 59800 2184
rect 200 1960 800 2156
rect 59200 1960 59800 2156
rect 130 1596 140 1652
rect 196 1596 2492 1652
rect 2548 1596 2558 1652
rect 200 1288 800 1512
rect 59200 1288 59800 1512
rect 200 616 800 840
rect 59200 616 59800 840
rect 58146 140 58156 196
rect 58212 168 59304 196
rect 58212 140 59800 168
rect 59200 -56 59800 140
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 52780 50428 52836 50484
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 52780 48636 52836 48692
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 52780 50484 52836 50494
rect 52780 48692 52836 50428
rect 52780 48626 52836 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__A1 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 56672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__A2
timestamp 1669390400
transform 1 0 56560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__A3
timestamp 1669390400
transform 1 0 53312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__A4
timestamp 1669390400
transform 1 0 57344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__A1
timestamp 1669390400
transform 1 0 55888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__A2
timestamp 1669390400
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__B1
timestamp 1669390400
transform 1 0 54544 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__B2
timestamp 1669390400
transform 1 0 54208 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__A1
timestamp 1669390400
transform -1 0 54432 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__A2
timestamp 1669390400
transform 1 0 53424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__A1
timestamp 1669390400
transform 1 0 53760 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A1
timestamp 1669390400
transform 1 0 54096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A2
timestamp 1669390400
transform 1 0 50960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A3
timestamp 1669390400
transform 1 0 50288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A1
timestamp 1669390400
transform -1 0 52640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A2
timestamp 1669390400
transform 1 0 50848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__B1
timestamp 1669390400
transform -1 0 51408 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__B2
timestamp 1669390400
transform -1 0 53088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A1
timestamp 1669390400
transform 1 0 50288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A2
timestamp 1669390400
transform 1 0 50736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__A1
timestamp 1669390400
transform 1 0 51632 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__A2
timestamp 1669390400
transform -1 0 52304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__A1
timestamp 1669390400
transform 1 0 54432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__A2
timestamp 1669390400
transform 1 0 53648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__A1
timestamp 1669390400
transform -1 0 49616 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__A2
timestamp 1669390400
transform 1 0 50624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A1
timestamp 1669390400
transform 1 0 51072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A2
timestamp 1669390400
transform 1 0 53312 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__B1
timestamp 1669390400
transform 1 0 52752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__B2
timestamp 1669390400
transform 1 0 54880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__A1
timestamp 1669390400
transform -1 0 53984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__A1
timestamp 1669390400
transform -1 0 53536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__A1
timestamp 1669390400
transform 1 0 54208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I
timestamp 1669390400
transform 1 0 53088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1669390400
transform 1 0 51744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__A1
timestamp 1669390400
transform 1 0 53536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__A1
timestamp 1669390400
transform 1 0 48384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__A2
timestamp 1669390400
transform 1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A1
timestamp 1669390400
transform 1 0 50288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A2
timestamp 1669390400
transform 1 0 50176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A3
timestamp 1669390400
transform 1 0 51520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A4
timestamp 1669390400
transform 1 0 50400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__A1
timestamp 1669390400
transform 1 0 50848 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__A2
timestamp 1669390400
transform 1 0 50848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__B1
timestamp 1669390400
transform 1 0 51296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__B2
timestamp 1669390400
transform 1 0 50400 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__A1
timestamp 1669390400
transform 1 0 49392 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__A2
timestamp 1669390400
transform 1 0 49728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__B1
timestamp 1669390400
transform 1 0 46928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__B2
timestamp 1669390400
transform 1 0 50176 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__A1
timestamp 1669390400
transform 1 0 51408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__A2
timestamp 1669390400
transform 1 0 47040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__C
timestamp 1669390400
transform 1 0 50736 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__A1
timestamp 1669390400
transform 1 0 50064 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__A2
timestamp 1669390400
transform 1 0 49616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__A3
timestamp 1669390400
transform 1 0 49168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__A1
timestamp 1669390400
transform 1 0 49280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__A2
timestamp 1669390400
transform 1 0 48720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__A1
timestamp 1669390400
transform 1 0 49168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__A2
timestamp 1669390400
transform -1 0 47040 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A1
timestamp 1669390400
transform -1 0 46256 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A2
timestamp 1669390400
transform 1 0 46480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__A1
timestamp 1669390400
transform -1 0 51408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__A2
timestamp 1669390400
transform 1 0 50848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__A1
timestamp 1669390400
transform -1 0 47488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__A2
timestamp 1669390400
transform 1 0 46256 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__A1
timestamp 1669390400
transform 1 0 45024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__I
timestamp 1669390400
transform -1 0 42896 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__A1
timestamp 1669390400
transform -1 0 44128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__A1
timestamp 1669390400
transform 1 0 49392 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__A2
timestamp 1669390400
transform 1 0 49392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__A1
timestamp 1669390400
transform 1 0 49392 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__A2
timestamp 1669390400
transform 1 0 48608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A1
timestamp 1669390400
transform -1 0 49728 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A2
timestamp 1669390400
transform -1 0 50176 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__A1
timestamp 1669390400
transform 1 0 50288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__A2
timestamp 1669390400
transform 1 0 49840 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__A1
timestamp 1669390400
transform 1 0 50624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__A2
timestamp 1669390400
transform 1 0 50176 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1669390400
transform -1 0 53648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A1
timestamp 1669390400
transform 1 0 44688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A2
timestamp 1669390400
transform 1 0 44016 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__A1
timestamp 1669390400
transform -1 0 44128 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__A2
timestamp 1669390400
transform 1 0 46368 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A1
timestamp 1669390400
transform 1 0 49840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A2
timestamp 1669390400
transform 1 0 49840 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1669390400
transform 1 0 56784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1669390400
transform 1 0 57344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1669390400
transform 1 0 50512 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__D
timestamp 1669390400
transform -1 0 46816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1669390400
transform 1 0 58016 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1669390400
transform 1 0 43568 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__D
timestamp 1669390400
transform 1 0 39424 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1669390400
transform 1 0 57568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__D
timestamp 1669390400
transform 1 0 58016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1669390400
transform 1 0 48832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1669390400
transform 1 0 56784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1669390400
transform 1 0 54544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__D
timestamp 1669390400
transform -1 0 54320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1669390400
transform 1 0 44912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__D
timestamp 1669390400
transform -1 0 40992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1669390400
transform 1 0 43232 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1669390400
transform -1 0 54768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1669390400
transform 1 0 53424 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1669390400
transform 1 0 50848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1669390400
transform 1 0 54768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1669390400
transform -1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1669390400
transform 1 0 42896 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1669390400
transform 1 0 54544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1669390400
transform -1 0 56336 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1669390400
transform 1 0 44912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout22_I
timestamp 1669390400
transform -1 0 55664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout23_I
timestamp 1669390400
transform 1 0 56784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout24_I
timestamp 1669390400
transform -1 0 55888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform 1 0 57344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 57568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 5824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 54096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform 1 0 57344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 45584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 56784 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform 1 0 57344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform 1 0 12992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform 1 0 57344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output12_I
timestamp 1669390400
transform 1 0 3472 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1669390400
transform 1 0 3696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1669390400
transform 1 0 50736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1669390400
transform -1 0 3696 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1669390400
transform 1 0 4816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1669390400
transform -1 0 15120 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17
timestamp 1669390400
transform 1 0 3248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23
timestamp 1669390400
transform 1 0 3920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29
timestamp 1669390400
transform 1 0 4592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33
timestamp 1669390400
transform 1 0 5040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_112 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120
timestamp 1669390400
transform 1 0 14784 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_125
timestamp 1669390400
transform 1 0 15344 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_137
timestamp 1669390400
transform 1 0 16688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_150
timestamp 1669390400
transform 1 0 18144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_154
timestamp 1669390400
transform 1 0 18592 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_156
timestamp 1669390400
transform 1 0 18816 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_161
timestamp 1669390400
transform 1 0 19376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169
timestamp 1669390400
transform 1 0 20272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1669390400
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_185
timestamp 1669390400
transform 1 0 22064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_191
timestamp 1669390400
transform 1 0 22736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_197
timestamp 1669390400
transform 1 0 23408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_228
timestamp 1669390400
transform 1 0 26880 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_236
timestamp 1669390400
transform 1 0 27776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1669390400
transform 1 0 28224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_264
timestamp 1669390400
transform 1 0 30912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_287
timestamp 1669390400
transform 1 0 33488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_295
timestamp 1669390400
transform 1 0 34384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_299
timestamp 1669390400
transform 1 0 34832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_305
timestamp 1669390400
transform 1 0 35504 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1669390400
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_322
timestamp 1669390400
transform 1 0 37408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_330
timestamp 1669390400
transform 1 0 38304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_334
timestamp 1669390400
transform 1 0 38752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_336
timestamp 1669390400
transform 1 0 38976 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_341
timestamp 1669390400
transform 1 0 39536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_347
timestamp 1669390400
transform 1 0 40208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_407
timestamp 1669390400
transform 1 0 46928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_413
timestamp 1669390400
transform 1 0 47600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1669390400
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_426
timestamp 1669390400
transform 1 0 49056 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_441
timestamp 1669390400
transform 1 0 50736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_447
timestamp 1669390400
transform 1 0 51408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1669390400
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_473
timestamp 1669390400
transform 1 0 54320 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_481
timestamp 1669390400
transform 1 0 55216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_497
timestamp 1669390400
transform 1 0 57008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_501
timestamp 1669390400
transform 1 0 57456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_503
timestamp 1669390400
transform 1 0 57680 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_508
timestamp 1669390400
transform 1 0 58240 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_7 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2128 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_89
timestamp 1669390400
transform 1 0 11312 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_101
timestamp 1669390400
transform 1 0 12656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_103
timestamp 1669390400
transform 1 0 12880 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_106
timestamp 1669390400
transform 1 0 13216 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_138
timestamp 1669390400
transform 1 0 16800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1669390400
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1669390400
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_436
timestamp 1669390400
transform 1 0 50176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_440
timestamp 1669390400
transform 1 0 50624 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_443
timestamp 1669390400
transform 1 0 50960 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_475
timestamp 1669390400
transform 1 0 54544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_493
timestamp 1669390400
transform 1 0 56560 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_502
timestamp 1669390400
transform 1 0 57568 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_508
timestamp 1669390400
transform 1 0 58240 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_7
timestamp 1669390400
transform 1 0 2128 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_23
timestamp 1669390400
transform 1 0 3920 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_31
timestamp 1669390400
transform 1 0 4816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1669390400
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1669390400
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_495
timestamp 1669390400
transform 1 0 56784 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_503
timestamp 1669390400
transform 1 0 57680 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_508
timestamp 1669390400
transform 1 0 58240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_503
timestamp 1669390400
transform 1 0 57680 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_508
timestamp 1669390400
transform 1 0 58240 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_7
timestamp 1669390400
transform 1 0 2128 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_23
timestamp 1669390400
transform 1 0 3920 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_31
timestamp 1669390400
transform 1 0 4816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_495
timestamp 1669390400
transform 1 0 56784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_503
timestamp 1669390400
transform 1 0 57680 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_507
timestamp 1669390400
transform 1 0 58128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_507
timestamp 1669390400
transform 1 0 58128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_495
timestamp 1669390400
transform 1 0 56784 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_503
timestamp 1669390400
transform 1 0 57680 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_507
timestamp 1669390400
transform 1 0 58128 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_507
timestamp 1669390400
transform 1 0 58128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_7
timestamp 1669390400
transform 1 0 2128 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_23
timestamp 1669390400
transform 1 0 3920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_31
timestamp 1669390400
transform 1 0 4816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_495
timestamp 1669390400
transform 1 0 56784 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_503
timestamp 1669390400
transform 1 0 57680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_507
timestamp 1669390400
transform 1 0 58128 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_7
timestamp 1669390400
transform 1 0 2128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_507
timestamp 1669390400
transform 1 0 58128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_495
timestamp 1669390400
transform 1 0 56784 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_503
timestamp 1669390400
transform 1 0 57680 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_508
timestamp 1669390400
transform 1 0 58240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_507
timestamp 1669390400
transform 1 0 58128 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_7
timestamp 1669390400
transform 1 0 2128 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_23
timestamp 1669390400
transform 1 0 3920 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_31
timestamp 1669390400
transform 1 0 4816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_495
timestamp 1669390400
transform 1 0 56784 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_503
timestamp 1669390400
transform 1 0 57680 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_507
timestamp 1669390400
transform 1 0 58128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_503
timestamp 1669390400
transform 1 0 57680 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_508
timestamp 1669390400
transform 1 0 58240 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_7
timestamp 1669390400
transform 1 0 2128 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_23
timestamp 1669390400
transform 1 0 3920 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_31
timestamp 1669390400
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_495
timestamp 1669390400
transform 1 0 56784 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_503
timestamp 1669390400
transform 1 0 57680 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_507
timestamp 1669390400
transform 1 0 58128 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_7
timestamp 1669390400
transform 1 0 2128 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_507
timestamp 1669390400
transform 1 0 58128 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_495
timestamp 1669390400
transform 1 0 56784 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_503
timestamp 1669390400
transform 1 0 57680 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_508
timestamp 1669390400
transform 1 0 58240 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_7
timestamp 1669390400
transform 1 0 2128 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_507
timestamp 1669390400
transform 1 0 58128 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_495
timestamp 1669390400
transform 1 0 56784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_503
timestamp 1669390400
transform 1 0 57680 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_507
timestamp 1669390400
transform 1 0 58128 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_7
timestamp 1669390400
transform 1 0 2128 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_507
timestamp 1669390400
transform 1 0 58128 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_495
timestamp 1669390400
transform 1 0 56784 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_503
timestamp 1669390400
transform 1 0 57680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_507
timestamp 1669390400
transform 1 0 58128 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_7
timestamp 1669390400
transform 1 0 2128 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_460
timestamp 1669390400
transform 1 0 52864 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_476
timestamp 1669390400
transform 1 0 54656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_493
timestamp 1669390400
transform 1 0 56560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_502
timestamp 1669390400
transform 1 0 57568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_506
timestamp 1669390400
transform 1 0 58016 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_508
timestamp 1669390400
transform 1 0 58240 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_495
timestamp 1669390400
transform 1 0 56784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_503
timestamp 1669390400
transform 1 0 57680 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_507
timestamp 1669390400
transform 1 0 58128 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_7
timestamp 1669390400
transform 1 0 2128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_507
timestamp 1669390400
transform 1 0 58128 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_7
timestamp 1669390400
transform 1 0 2128 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_23
timestamp 1669390400
transform 1 0 3920 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_31
timestamp 1669390400
transform 1 0 4816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_495
timestamp 1669390400
transform 1 0 56784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_503
timestamp 1669390400
transform 1 0 57680 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_507
timestamp 1669390400
transform 1 0 58128 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_7
timestamp 1669390400
transform 1 0 2128 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_460
timestamp 1669390400
transform 1 0 52864 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_476
timestamp 1669390400
transform 1 0 54656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_493
timestamp 1669390400
transform 1 0 56560 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_502
timestamp 1669390400
transform 1 0 57568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_506
timestamp 1669390400
transform 1 0 58016 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_508
timestamp 1669390400
transform 1 0 58240 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_495
timestamp 1669390400
transform 1 0 56784 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_503
timestamp 1669390400
transform 1 0 57680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_507
timestamp 1669390400
transform 1 0 58128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_503
timestamp 1669390400
transform 1 0 57680 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_508
timestamp 1669390400
transform 1 0 58240 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_17
timestamp 1669390400
transform 1 0 3248 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_21
timestamp 1669390400
transform 1 0 3696 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_29
timestamp 1669390400
transform 1 0 4592 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_33
timestamp 1669390400
transform 1 0 5040 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_337
timestamp 1669390400
transform 1 0 39088 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_345
timestamp 1669390400
transform 1 0 39984 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_347
timestamp 1669390400
transform 1 0 40208 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_377
timestamp 1669390400
transform 1 0 43568 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_381
timestamp 1669390400
transform 1 0 44016 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_495
timestamp 1669390400
transform 1 0 56784 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_503
timestamp 1669390400
transform 1 0 57680 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_507
timestamp 1669390400
transform 1 0 58128 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_367
timestamp 1669390400
transform 1 0 42448 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_371
timestamp 1669390400
transform 1 0 42896 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_403
timestamp 1669390400
transform 1 0 46480 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_419
timestamp 1669390400
transform 1 0 48272 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_423
timestamp 1669390400
transform 1 0 48720 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_507
timestamp 1669390400
transform 1 0 58128 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_7
timestamp 1669390400
transform 1 0 2128 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_23
timestamp 1669390400
transform 1 0 3920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_31
timestamp 1669390400
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_495
timestamp 1669390400
transform 1 0 56784 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_503
timestamp 1669390400
transform 1 0 57680 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_507
timestamp 1669390400
transform 1 0 58128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_507
timestamp 1669390400
transform 1 0 58128 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_7
timestamp 1669390400
transform 1 0 2128 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_23
timestamp 1669390400
transform 1 0 3920 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_31
timestamp 1669390400
transform 1 0 4816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_495
timestamp 1669390400
transform 1 0 56784 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_503
timestamp 1669390400
transform 1 0 57680 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_508
timestamp 1669390400
transform 1 0 58240 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_507
timestamp 1669390400
transform 1 0 58128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_495
timestamp 1669390400
transform 1 0 56784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_503
timestamp 1669390400
transform 1 0 57680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_507
timestamp 1669390400
transform 1 0 58128 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_503
timestamp 1669390400
transform 1 0 57680 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_508
timestamp 1669390400
transform 1 0 58240 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_7
timestamp 1669390400
transform 1 0 2128 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_13
timestamp 1669390400
transform 1 0 2800 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_29
timestamp 1669390400
transform 1 0 4592 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_33
timestamp 1669390400
transform 1 0 5040 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_495
timestamp 1669390400
transform 1 0 56784 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_497
timestamp 1669390400
transform 1 0 57008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_502
timestamp 1669390400
transform 1 0 57568 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_508
timestamp 1669390400
transform 1 0 58240 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_507
timestamp 1669390400
transform 1 0 58128 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_495
timestamp 1669390400
transform 1 0 56784 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_503
timestamp 1669390400
transform 1 0 57680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_507
timestamp 1669390400
transform 1 0 58128 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_507
timestamp 1669390400
transform 1 0 58128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_471
timestamp 1669390400
transform 1 0 54096 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_477
timestamp 1669390400
transform 1 0 54768 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_508
timestamp 1669390400
transform 1 0 58240 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_7
timestamp 1669390400
transform 1 0 2128 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_460
timestamp 1669390400
transform 1 0 52864 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_476
timestamp 1669390400
transform 1 0 54656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_491
timestamp 1669390400
transform 1 0 56336 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_495
timestamp 1669390400
transform 1 0 56784 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_507
timestamp 1669390400
transform 1 0 58128 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_408
timestamp 1669390400
transform 1 0 47040 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_410
timestamp 1669390400
transform 1 0 47264 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_440
timestamp 1669390400
transform 1 0 50624 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_444
timestamp 1669390400
transform 1 0 51072 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_471
timestamp 1669390400
transform 1 0 54096 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_475
timestamp 1669390400
transform 1 0 54544 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_483
timestamp 1669390400
transform 1 0 55440 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_487
timestamp 1669390400
transform 1 0 55888 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_503
timestamp 1669390400
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_507
timestamp 1669390400
transform 1 0 58128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_460
timestamp 1669390400
transform 1 0 52864 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_464
timestamp 1669390400
transform 1 0 53312 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_467
timestamp 1669390400
transform 1 0 53648 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_475
timestamp 1669390400
transform 1 0 54544 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_493
timestamp 1669390400
transform 1 0 56560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_502
timestamp 1669390400
transform 1 0 57568 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_506
timestamp 1669390400
transform 1 0 58016 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_508
timestamp 1669390400
transform 1 0 58240 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1669390400
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_493
timestamp 1669390400
transform 1 0 56560 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_497
timestamp 1669390400
transform 1 0 57008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_505
timestamp 1669390400
transform 1 0 57904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1669390400
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_435
timestamp 1669390400
transform 1 0 50064 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_439
timestamp 1669390400
transform 1 0 50512 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_469
timestamp 1669390400
transform 1 0 53872 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_473
timestamp 1669390400
transform 1 0 54320 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_477
timestamp 1669390400
transform 1 0 54768 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_493
timestamp 1669390400
transform 1 0 56560 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_507
timestamp 1669390400
transform 1 0 58128 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_7
timestamp 1669390400
transform 1 0 2128 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_23
timestamp 1669390400
transform 1 0 3920 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_31
timestamp 1669390400
transform 1 0 4816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1669390400
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_408
timestamp 1669390400
transform 1 0 47040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_412
timestamp 1669390400
transform 1 0 47488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_422
timestamp 1669390400
transform 1 0 48608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_426
timestamp 1669390400
transform 1 0 49056 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_440
timestamp 1669390400
transform 1 0 50624 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_444
timestamp 1669390400
transform 1 0 51072 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_495
timestamp 1669390400
transform 1 0 56784 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_503
timestamp 1669390400
transform 1 0 57680 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_508
timestamp 1669390400
transform 1 0 58240 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_7
timestamp 1669390400
transform 1 0 2128 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_350
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_387
timestamp 1669390400
transform 1 0 44688 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_391
timestamp 1669390400
transform 1 0 45136 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_399
timestamp 1669390400
transform 1 0 46032 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_403
timestamp 1669390400
transform 1 0 46480 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_410
timestamp 1669390400
transform 1 0 47264 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_414
timestamp 1669390400
transform 1 0 47712 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_420
timestamp 1669390400
transform 1 0 48384 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_424
timestamp 1669390400
transform 1 0 48832 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_435
timestamp 1669390400
transform 1 0 50064 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_439
timestamp 1669390400
transform 1 0 50512 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_443
timestamp 1669390400
transform 1 0 50960 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_447
timestamp 1669390400
transform 1 0 51408 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_451
timestamp 1669390400
transform 1 0 51856 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_455
timestamp 1669390400
transform 1 0 52304 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_471
timestamp 1669390400
transform 1 0 54096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_475
timestamp 1669390400
transform 1 0 54544 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_491
timestamp 1669390400
transform 1 0 56336 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_495
timestamp 1669390400
transform 1 0 56784 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_503
timestamp 1669390400
transform 1 0 57680 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_508
timestamp 1669390400
transform 1 0 58240 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_7
timestamp 1669390400
transform 1 0 2128 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_13
timestamp 1669390400
transform 1 0 2800 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_29
timestamp 1669390400
transform 1 0 4592 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_33
timestamp 1669390400
transform 1 0 5040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_394
timestamp 1669390400
transform 1 0 45472 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_407
timestamp 1669390400
transform 1 0 46928 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_414
timestamp 1669390400
transform 1 0 47712 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_427
timestamp 1669390400
transform 1 0 49168 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_434
timestamp 1669390400
transform 1 0 49952 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_438
timestamp 1669390400
transform 1 0 50400 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_440
timestamp 1669390400
transform 1 0 50624 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_446
timestamp 1669390400
transform 1 0 51296 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_450
timestamp 1669390400
transform 1 0 51744 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_466
timestamp 1669390400
transform 1 0 53536 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_470
timestamp 1669390400
transform 1 0 53984 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_474
timestamp 1669390400
transform 1 0 54432 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_477
timestamp 1669390400
transform 1 0 54768 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_508
timestamp 1669390400
transform 1 0 58240 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_389
timestamp 1669390400
transform 1 0 44912 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_393
timestamp 1669390400
transform 1 0 45360 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_395
timestamp 1669390400
transform 1 0 45584 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_408
timestamp 1669390400
transform 1 0 47040 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_412
timestamp 1669390400
transform 1 0 47488 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_435
timestamp 1669390400
transform 1 0 50064 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_439
timestamp 1669390400
transform 1 0 50512 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_464
timestamp 1669390400
transform 1 0 53312 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_481
timestamp 1669390400
transform 1 0 55216 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_507
timestamp 1669390400
transform 1 0 58128 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_337
timestamp 1669390400
transform 1 0 39088 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_339
timestamp 1669390400
transform 1 0 39312 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_342
timestamp 1669390400
transform 1 0 39648 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_375
timestamp 1669390400
transform 1 0 43344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_379
timestamp 1669390400
transform 1 0 43792 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_387
timestamp 1669390400
transform 1 0 44688 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_396
timestamp 1669390400
transform 1 0 45696 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_398
timestamp 1669390400
transform 1 0 45920 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_407
timestamp 1669390400
transform 1 0 46928 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_425
timestamp 1669390400
transform 1 0 48944 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_436
timestamp 1669390400
transform 1 0 50176 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_440
timestamp 1669390400
transform 1 0 50624 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_444
timestamp 1669390400
transform 1 0 51072 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_446
timestamp 1669390400
transform 1 0 51296 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_451
timestamp 1669390400
transform 1 0 51856 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_457
timestamp 1669390400
transform 1 0 52528 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_470
timestamp 1669390400
transform 1 0 53984 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_474
timestamp 1669390400
transform 1 0 54432 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_476
timestamp 1669390400
transform 1 0 54656 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_493
timestamp 1669390400
transform 1 0 56560 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_497
timestamp 1669390400
transform 1 0 57008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_505
timestamp 1669390400
transform 1 0 57904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_373
timestamp 1669390400
transform 1 0 43120 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_377
timestamp 1669390400
transform 1 0 43568 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_379
timestamp 1669390400
transform 1 0 43792 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_382
timestamp 1669390400
transform 1 0 44128 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_390
timestamp 1669390400
transform 1 0 45024 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_392
timestamp 1669390400
transform 1 0 45248 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_405
timestamp 1669390400
transform 1 0 46704 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_409
timestamp 1669390400
transform 1 0 47152 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_411
timestamp 1669390400
transform 1 0 47376 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_436
timestamp 1669390400
transform 1 0 50176 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_440
timestamp 1669390400
transform 1 0 50624 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_444
timestamp 1669390400
transform 1 0 51072 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_448
timestamp 1669390400
transform 1 0 51520 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_452
timestamp 1669390400
transform 1 0 51968 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_454
timestamp 1669390400
transform 1 0 52192 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_460
timestamp 1669390400
transform 1 0 52864 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_464
timestamp 1669390400
transform 1 0 53312 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_468
timestamp 1669390400
transform 1 0 53760 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_484
timestamp 1669390400
transform 1 0 55552 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1669390400
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_501
timestamp 1669390400
transform 1 0 57456 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_504
timestamp 1669390400
transform 1 0 57792 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_508
timestamp 1669390400
transform 1 0 58240 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_353
timestamp 1669390400
transform 1 0 40880 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_369
timestamp 1669390400
transform 1 0 42672 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_373
timestamp 1669390400
transform 1 0 43120 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_380
timestamp 1669390400
transform 1 0 43904 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_382
timestamp 1669390400
transform 1 0 44128 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_405
timestamp 1669390400
transform 1 0 46704 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_407
timestamp 1669390400
transform 1 0 46928 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_410
timestamp 1669390400
transform 1 0 47264 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_445
timestamp 1669390400
transform 1 0 51184 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_449
timestamp 1669390400
transform 1 0 51632 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_472
timestamp 1669390400
transform 1 0 54208 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_476
timestamp 1669390400
transform 1 0 54656 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_508
timestamp 1669390400
transform 1 0 58240 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_7
timestamp 1669390400
transform 1 0 2128 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_361
timestamp 1669390400
transform 1 0 41776 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_374
timestamp 1669390400
transform 1 0 43232 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_388
timestamp 1669390400
transform 1 0 44800 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_392
timestamp 1669390400
transform 1 0 45248 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_406
timestamp 1669390400
transform 1 0 46816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_410
timestamp 1669390400
transform 1 0 47264 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_431
timestamp 1669390400
transform 1 0 49616 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_439
timestamp 1669390400
transform 1 0 50512 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_443
timestamp 1669390400
transform 1 0 50960 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_457
timestamp 1669390400
transform 1 0 52528 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_483
timestamp 1669390400
transform 1 0 55440 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_493
timestamp 1669390400
transform 1 0 56560 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_503
timestamp 1669390400
transform 1 0 57680 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_508
timestamp 1669390400
transform 1 0 58240 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_7
timestamp 1669390400
transform 1 0 2128 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_13
timestamp 1669390400
transform 1 0 2800 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_29
timestamp 1669390400
transform 1 0 4592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_33
timestamp 1669390400
transform 1 0 5040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1669390400
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1669390400
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_353
timestamp 1669390400
transform 1 0 40880 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_377
timestamp 1669390400
transform 1 0 43568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1669390400
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1669390400
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_396
timestamp 1669390400
transform 1 0 45696 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_398
timestamp 1669390400
transform 1 0 45920 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_403
timestamp 1669390400
transform 1 0 46480 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_407
timestamp 1669390400
transform 1 0 46928 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_412
timestamp 1669390400
transform 1 0 47488 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_425
timestamp 1669390400
transform 1 0 48944 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_429
timestamp 1669390400
transform 1 0 49392 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_433
timestamp 1669390400
transform 1 0 49840 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_437
timestamp 1669390400
transform 1 0 50288 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_439
timestamp 1669390400
transform 1 0 50512 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_448
timestamp 1669390400
transform 1 0 51520 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_458
timestamp 1669390400
transform 1 0 52640 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_472
timestamp 1669390400
transform 1 0 54208 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_476
timestamp 1669390400
transform 1 0 54656 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_480
timestamp 1669390400
transform 1 0 55104 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_482
timestamp 1669390400
transform 1 0 55328 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_485
timestamp 1669390400
transform 1 0 55664 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_489
timestamp 1669390400
transform 1 0 56112 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_497
timestamp 1669390400
transform 1 0 57008 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_499
timestamp 1669390400
transform 1 0 57232 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_502
timestamp 1669390400
transform 1 0 57568 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_508
timestamp 1669390400
transform 1 0 58240 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1669390400
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1669390400
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1669390400
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1669390400
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_389
timestamp 1669390400
transform 1 0 44912 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_397
timestamp 1669390400
transform 1 0 45808 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_401
timestamp 1669390400
transform 1 0 46256 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_405
timestamp 1669390400
transform 1 0 46704 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_414
timestamp 1669390400
transform 1 0 47712 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_438
timestamp 1669390400
transform 1 0 50400 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_451
timestamp 1669390400
transform 1 0 51856 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_458
timestamp 1669390400
transform 1 0 52640 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_465
timestamp 1669390400
transform 1 0 53424 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_469
timestamp 1669390400
transform 1 0 53872 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_473
timestamp 1669390400
transform 1 0 54320 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_480
timestamp 1669390400
transform 1 0 55104 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_488
timestamp 1669390400
transform 1 0 56000 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_492
timestamp 1669390400
transform 1 0 56448 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_502
timestamp 1669390400
transform 1 0 57568 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_508
timestamp 1669390400
transform 1 0 58240 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_7
timestamp 1669390400
transform 1 0 2128 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_23
timestamp 1669390400
transform 1 0 3920 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_31
timestamp 1669390400
transform 1 0 4816 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1669390400
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_353
timestamp 1669390400
transform 1 0 40880 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_361
timestamp 1669390400
transform 1 0 41776 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_365
timestamp 1669390400
transform 1 0 42224 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_379
timestamp 1669390400
transform 1 0 43792 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_386
timestamp 1669390400
transform 1 0 44576 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_405
timestamp 1669390400
transform 1 0 46704 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_409
timestamp 1669390400
transform 1 0 47152 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_419
timestamp 1669390400
transform 1 0 48272 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_426
timestamp 1669390400
transform 1 0 49056 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_430
timestamp 1669390400
transform 1 0 49504 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_434
timestamp 1669390400
transform 1 0 49952 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_438
timestamp 1669390400
transform 1 0 50400 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_442
timestamp 1669390400
transform 1 0 50848 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_446
timestamp 1669390400
transform 1 0 51296 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_448
timestamp 1669390400
transform 1 0 51520 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_457
timestamp 1669390400
transform 1 0 52528 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_466
timestamp 1669390400
transform 1 0 53536 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_477
timestamp 1669390400
transform 1 0 54768 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_508
timestamp 1669390400
transform 1 0 58240 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1669390400
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1669390400
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_371
timestamp 1669390400
transform 1 0 42896 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_375
timestamp 1669390400
transform 1 0 43344 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_377
timestamp 1669390400
transform 1 0 43568 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_390
timestamp 1669390400
transform 1 0 45024 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_407
timestamp 1669390400
transform 1 0 46928 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_415
timestamp 1669390400
transform 1 0 47824 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_421
timestamp 1669390400
transform 1 0 48496 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_431
timestamp 1669390400
transform 1 0 49616 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_435
timestamp 1669390400
transform 1 0 50064 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_439
timestamp 1669390400
transform 1 0 50512 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_445
timestamp 1669390400
transform 1 0 51184 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_457
timestamp 1669390400
transform 1 0 52528 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_461
timestamp 1669390400
transform 1 0 52976 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_463
timestamp 1669390400
transform 1 0 53200 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_475
timestamp 1669390400
transform 1 0 54544 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_493
timestamp 1669390400
transform 1 0 56560 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_502
timestamp 1669390400
transform 1 0 57568 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_508
timestamp 1669390400
transform 1 0 58240 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1669390400
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1669390400
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_359
timestamp 1669390400
transform 1 0 41552 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_375
timestamp 1669390400
transform 1 0 43344 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_404
timestamp 1669390400
transform 1 0 46592 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_408
timestamp 1669390400
transform 1 0 47040 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_415
timestamp 1669390400
transform 1 0 47824 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_425
timestamp 1669390400
transform 1 0 48944 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_429
timestamp 1669390400
transform 1 0 49392 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_433
timestamp 1669390400
transform 1 0 49840 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_445
timestamp 1669390400
transform 1 0 51184 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_469
timestamp 1669390400
transform 1 0 53872 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_473
timestamp 1669390400
transform 1 0 54320 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_477
timestamp 1669390400
transform 1 0 54768 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_508
timestamp 1669390400
transform 1 0 58240 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_373
timestamp 1669390400
transform 1 0 43120 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_381
timestamp 1669390400
transform 1 0 44016 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_391
timestamp 1669390400
transform 1 0 45136 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_399
timestamp 1669390400
transform 1 0 46032 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_407
timestamp 1669390400
transform 1 0 46928 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_418
timestamp 1669390400
transform 1 0 48160 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_431
timestamp 1669390400
transform 1 0 49616 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_435
timestamp 1669390400
transform 1 0 50064 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_445
timestamp 1669390400
transform 1 0 51184 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_456
timestamp 1669390400
transform 1 0 52416 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_463
timestamp 1669390400
transform 1 0 53200 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_470
timestamp 1669390400
transform 1 0 53984 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_474
timestamp 1669390400
transform 1 0 54432 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_476
timestamp 1669390400
transform 1 0 54656 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_491
timestamp 1669390400
transform 1 0 56336 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_495
timestamp 1669390400
transform 1 0 56784 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_503
timestamp 1669390400
transform 1 0 57680 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_505
timestamp 1669390400
transform 1 0 57904 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_508
timestamp 1669390400
transform 1 0 58240 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1669390400
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_337
timestamp 1669390400
transform 1 0 39088 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_339
timestamp 1669390400
transform 1 0 39312 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_369
timestamp 1669390400
transform 1 0 42672 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_373
timestamp 1669390400
transform 1 0 43120 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_381
timestamp 1669390400
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_385
timestamp 1669390400
transform 1 0 44464 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_406
timestamp 1669390400
transform 1 0 46816 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_420
timestamp 1669390400
transform 1 0 48384 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_427
timestamp 1669390400
transform 1 0 49168 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_431
timestamp 1669390400
transform 1 0 49616 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_435
timestamp 1669390400
transform 1 0 50064 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_439
timestamp 1669390400
transform 1 0 50512 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_441
timestamp 1669390400
transform 1 0 50736 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_444
timestamp 1669390400
transform 1 0 51072 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_459
timestamp 1669390400
transform 1 0 52752 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_466
timestamp 1669390400
transform 1 0 53536 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_470
timestamp 1669390400
transform 1 0 53984 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_474
timestamp 1669390400
transform 1 0 54432 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_478
timestamp 1669390400
transform 1 0 54880 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_508
timestamp 1669390400
transform 1 0 58240 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_7
timestamp 1669390400
transform 1 0 2128 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1669390400
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_364
timestamp 1669390400
transform 1 0 42112 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_380
timestamp 1669390400
transform 1 0 43904 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_383
timestamp 1669390400
transform 1 0 44240 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_390
timestamp 1669390400
transform 1 0 45024 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_394
timestamp 1669390400
transform 1 0 45472 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_400
timestamp 1669390400
transform 1 0 46144 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_407
timestamp 1669390400
transform 1 0 46928 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_422
timestamp 1669390400
transform 1 0 48608 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_434
timestamp 1669390400
transform 1 0 49952 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_438
timestamp 1669390400
transform 1 0 50400 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_442
timestamp 1669390400
transform 1 0 50848 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_444
timestamp 1669390400
transform 1 0 51072 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_447
timestamp 1669390400
transform 1 0 51408 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_455
timestamp 1669390400
transform 1 0 52304 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_458
timestamp 1669390400
transform 1 0 52640 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_462
timestamp 1669390400
transform 1 0 53088 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_464
timestamp 1669390400
transform 1 0 53312 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_467
timestamp 1669390400
transform 1 0 53648 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_475
timestamp 1669390400
transform 1 0 54544 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_479
timestamp 1669390400
transform 1 0 54992 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_495
timestamp 1669390400
transform 1 0 56784 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_503
timestamp 1669390400
transform 1 0 57680 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_508
timestamp 1669390400
transform 1 0 58240 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_337
timestamp 1669390400
transform 1 0 39088 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_341
timestamp 1669390400
transform 1 0 39536 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_372
timestamp 1669390400
transform 1 0 43008 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_376
timestamp 1669390400
transform 1 0 43456 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_382
timestamp 1669390400
transform 1 0 44128 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_400
timestamp 1669390400
transform 1 0 46144 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_404
timestamp 1669390400
transform 1 0 46592 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_408
timestamp 1669390400
transform 1 0 47040 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_421
timestamp 1669390400
transform 1 0 48496 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_428
timestamp 1669390400
transform 1 0 49280 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_432
timestamp 1669390400
transform 1 0 49728 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_436
timestamp 1669390400
transform 1 0 50176 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_444
timestamp 1669390400
transform 1 0 51072 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_451
timestamp 1669390400
transform 1 0 51856 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_459
timestamp 1669390400
transform 1 0 52752 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_493
timestamp 1669390400
transform 1 0 56560 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_497
timestamp 1669390400
transform 1 0 57008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_505
timestamp 1669390400
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_7
timestamp 1669390400
transform 1 0 2128 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_373
timestamp 1669390400
transform 1 0 43120 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_389
timestamp 1669390400
transform 1 0 44912 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_391
timestamp 1669390400
transform 1 0 45136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_397
timestamp 1669390400
transform 1 0 45808 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_413
timestamp 1669390400
transform 1 0 47600 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_420
timestamp 1669390400
transform 1 0 48384 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_424
timestamp 1669390400
transform 1 0 48832 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_431
timestamp 1669390400
transform 1 0 49616 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_433
timestamp 1669390400
transform 1 0 49840 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_463
timestamp 1669390400
transform 1 0 53200 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_467
timestamp 1669390400
transform 1 0 53648 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_483
timestamp 1669390400
transform 1 0 55440 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_491
timestamp 1669390400
transform 1 0 56336 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_495
timestamp 1669390400
transform 1 0 56784 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_503
timestamp 1669390400
transform 1 0 57680 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_508
timestamp 1669390400
transform 1 0 58240 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_17
timestamp 1669390400
transform 1 0 3248 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_21
timestamp 1669390400
transform 1 0 3696 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_29
timestamp 1669390400
transform 1 0 4592 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_33
timestamp 1669390400
transform 1 0 5040 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_353
timestamp 1669390400
transform 1 0 40880 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_369
timestamp 1669390400
transform 1 0 42672 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_400
timestamp 1669390400
transform 1 0 46144 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_406
timestamp 1669390400
transform 1 0 46816 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_437
timestamp 1669390400
transform 1 0 50288 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_441
timestamp 1669390400
transform 1 0 50736 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_457
timestamp 1669390400
transform 1 0 52528 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_495
timestamp 1669390400
transform 1 0 56784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_503
timestamp 1669390400
transform 1 0 57680 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_508
timestamp 1669390400
transform 1 0 58240 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_7
timestamp 1669390400
transform 1 0 2128 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_13
timestamp 1669390400
transform 1 0 2800 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_19
timestamp 1669390400
transform 1 0 3472 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_23
timestamp 1669390400
transform 1 0 3920 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_55
timestamp 1669390400
transform 1 0 7504 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_387
timestamp 1669390400
transform 1 0 44688 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_391
timestamp 1669390400
transform 1 0 45136 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_423
timestamp 1669390400
transform 1 0 48720 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_444
timestamp 1669390400
transform 1 0 51072 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_448
timestamp 1669390400
transform 1 0 51520 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_456
timestamp 1669390400
transform 1 0 52416 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_487
timestamp 1669390400
transform 1 0 55888 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_491
timestamp 1669390400
transform 1 0 56336 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_495
timestamp 1669390400
transform 1 0 56784 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_503
timestamp 1669390400
transform 1 0 57680 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_508
timestamp 1669390400
transform 1 0 58240 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_17
timestamp 1669390400
transform 1 0 3248 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_23
timestamp 1669390400
transform 1 0 3920 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_29
timestamp 1669390400
transform 1 0 4592 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_33
timestamp 1669390400
transform 1 0 5040 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_40
timestamp 1669390400
transform 1 0 5824 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_104
timestamp 1669390400
transform 1 0 12992 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_113
timestamp 1669390400
transform 1 0 14000 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1669390400
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1669390400
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1669390400
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_422
timestamp 1669390400
transform 1 0 48608 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_426
timestamp 1669390400
transform 1 0 49056 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_458
timestamp 1669390400
transform 1 0 52640 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1669390400
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_471
timestamp 1669390400
transform 1 0 54096 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_475
timestamp 1669390400
transform 1 0 54544 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_493
timestamp 1669390400
transform 1 0 56560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_497
timestamp 1669390400
transform 1 0 57008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_502
timestamp 1669390400
transform 1 0 57568 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_508
timestamp 1669390400
transform 1 0 58240 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_7
timestamp 1669390400
transform 1 0 2128 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_11
timestamp 1669390400
transform 1 0 2576 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_27
timestamp 1669390400
transform 1 0 4368 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_29
timestamp 1669390400
transform 1 0 4592 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_34
timestamp 1669390400
transform 1 0 5152 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_37
timestamp 1669390400
transform 1 0 5488 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_54
timestamp 1669390400
transform 1 0 7392 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_72
timestamp 1669390400
transform 1 0 9408 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_77
timestamp 1669390400
transform 1 0 9968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_81
timestamp 1669390400
transform 1 0 10416 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_83
timestamp 1669390400
transform 1 0 10640 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_88
timestamp 1669390400
transform 1 0 11200 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_104
timestamp 1669390400
transform 1 0 12992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_107
timestamp 1669390400
transform 1 0 13328 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_113
timestamp 1669390400
transform 1 0 14000 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_119
timestamp 1669390400
transform 1 0 14672 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_123
timestamp 1669390400
transform 1 0 15120 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_131
timestamp 1669390400
transform 1 0 16016 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1669390400
transform 1 0 16912 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_142
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_150
timestamp 1669390400
transform 1 0 18144 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_154
timestamp 1669390400
transform 1 0 18592 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_156
timestamp 1669390400
transform 1 0 18816 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_161
timestamp 1669390400
transform 1 0 19376 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_167
timestamp 1669390400
transform 1 0 20048 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_177
timestamp 1669390400
transform 1 0 21168 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_182
timestamp 1669390400
transform 1 0 21728 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_186
timestamp 1669390400
transform 1 0 22176 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_191
timestamp 1669390400
transform 1 0 22736 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_207
timestamp 1669390400
transform 1 0 24528 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_209
timestamp 1669390400
transform 1 0 24752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_228
timestamp 1669390400
transform 1 0 26880 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_233
timestamp 1669390400
transform 1 0 27440 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_237
timestamp 1669390400
transform 1 0 27888 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_239
timestamp 1669390400
transform 1 0 28112 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_244
timestamp 1669390400
transform 1 0 28672 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_247
timestamp 1669390400
transform 1 0 29008 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_251
timestamp 1669390400
transform 1 0 29456 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_257
timestamp 1669390400
transform 1 0 30128 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_265
timestamp 1669390400
transform 1 0 31024 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_269
timestamp 1669390400
transform 1 0 31472 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_275
timestamp 1669390400
transform 1 0 32144 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_282
timestamp 1669390400
transform 1 0 32928 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_287
timestamp 1669390400
transform 1 0 33488 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_293
timestamp 1669390400
transform 1 0 34160 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_309
timestamp 1669390400
transform 1 0 35952 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_313
timestamp 1669390400
transform 1 0 36400 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_317
timestamp 1669390400
transform 1 0 36848 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_322
timestamp 1669390400
transform 1 0 37408 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_328
timestamp 1669390400
transform 1 0 38080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_330
timestamp 1669390400
transform 1 0 38304 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_335
timestamp 1669390400
transform 1 0 38864 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_341
timestamp 1669390400
transform 1 0 39536 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_349
timestamp 1669390400
transform 1 0 40432 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_352
timestamp 1669390400
transform 1 0 40768 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_363
timestamp 1669390400
transform 1 0 42000 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_383
timestamp 1669390400
transform 1 0 44240 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_387
timestamp 1669390400
transform 1 0 44688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_391
timestamp 1669390400
transform 1 0 45136 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_395
timestamp 1669390400
transform 1 0 45584 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_413
timestamp 1669390400
transform 1 0 47600 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_419
timestamp 1669390400
transform 1 0 48272 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_422
timestamp 1669390400
transform 1 0 48608 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_427
timestamp 1669390400
transform 1 0 49168 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_433
timestamp 1669390400
transform 1 0 49840 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_449
timestamp 1669390400
transform 1 0 51632 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_453
timestamp 1669390400
transform 1 0 52080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_457
timestamp 1669390400
transform 1 0 52528 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_465
timestamp 1669390400
transform 1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_471
timestamp 1669390400
transform 1 0 54096 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_489
timestamp 1669390400
transform 1 0 56112 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_507
timestamp 1669390400
transform 1 0 58128 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 5264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 28784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 44464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 52304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _095_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53312 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _096_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53760 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _097_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54432 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _098_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 53200 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 50288 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _100_
timestamp 1669390400
transform -1 0 53872 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _101_
timestamp 1669390400
transform 1 0 49952 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _102_
timestamp 1669390400
transform 1 0 51408 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _103_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51408 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _104_
timestamp 1669390400
transform -1 0 53984 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _105_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 52752 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51184 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _107_
timestamp 1669390400
transform 1 0 49504 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _108_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51408 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _109_
timestamp 1669390400
transform -1 0 51296 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _110_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51632 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _111_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 50624 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _112_
timestamp 1669390400
transform -1 0 50400 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _113_
timestamp 1669390400
transform 1 0 50848 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _114_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51744 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _115_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51184 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _116_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 50736 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _117_
timestamp 1669390400
transform -1 0 50624 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1669390400
transform -1 0 50064 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _119_
timestamp 1669390400
transform 1 0 51968 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _120_
timestamp 1669390400
transform 1 0 53312 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _121_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 52080 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _122_
timestamp 1669390400
transform 1 0 51408 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  _123_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53536 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1669390400
transform 1 0 52080 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1669390400
transform -1 0 52864 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1669390400
transform 1 0 52864 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1669390400
transform 1 0 47824 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _128_
timestamp 1669390400
transform 1 0 47936 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _129_
timestamp 1669390400
transform -1 0 50176 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _130_
timestamp 1669390400
transform -1 0 50064 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _131_
timestamp 1669390400
transform -1 0 48944 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _132_
timestamp 1669390400
transform -1 0 48944 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _133_
timestamp 1669390400
transform 1 0 47040 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _134_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 51184 0 1 43904
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _135_
timestamp 1669390400
transform -1 0 48944 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _136_
timestamp 1669390400
transform 1 0 47488 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _137_
timestamp 1669390400
transform 1 0 47488 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _138_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 52752 0 -1 45472
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _139_
timestamp 1669390400
transform 1 0 55328 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _140_
timestamp 1669390400
transform -1 0 49056 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1669390400
transform 1 0 47264 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _142_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 47712 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1669390400
transform -1 0 48496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _144_
timestamp 1669390400
transform 1 0 47376 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _145_
timestamp 1669390400
transform 1 0 52080 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _146_
timestamp 1669390400
transform 1 0 53312 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_
timestamp 1669390400
transform 1 0 53312 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _148_
timestamp 1669390400
transform -1 0 44912 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _149_
timestamp 1669390400
transform -1 0 49952 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _150_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 48944 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1669390400
transform -1 0 47264 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _152_
timestamp 1669390400
transform 1 0 45696 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _153_
timestamp 1669390400
transform -1 0 46928 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _154_
timestamp 1669390400
transform -1 0 46704 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _155_
timestamp 1669390400
transform -1 0 46704 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _156_
timestamp 1669390400
transform -1 0 44800 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _157_
timestamp 1669390400
transform -1 0 43232 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _158_
timestamp 1669390400
transform 1 0 41776 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _159_
timestamp 1669390400
transform -1 0 43904 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _160_
timestamp 1669390400
transform 1 0 42672 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1669390400
transform 1 0 46032 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _162_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 45472 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1669390400
transform 1 0 47152 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 46032 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1669390400
transform -1 0 48944 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1669390400
transform -1 0 48384 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1669390400
transform -1 0 49280 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _168_
timestamp 1669390400
transform -1 0 48608 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _169_
timestamp 1669390400
transform -1 0 48384 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _170_
timestamp 1669390400
transform 1 0 45472 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _171_
timestamp 1669390400
transform -1 0 46704 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _172_
timestamp 1669390400
transform -1 0 43792 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _173_
timestamp 1669390400
transform -1 0 42896 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _174_
timestamp 1669390400
transform 1 0 40880 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1669390400
transform -1 0 44576 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _176_
timestamp 1669390400
transform 1 0 42448 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _177_
timestamp 1669390400
transform 1 0 47152 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _178_
timestamp 1669390400
transform 1 0 45696 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _179_
timestamp 1669390400
transform -1 0 49168 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _180_
timestamp 1669390400
transform -1 0 48160 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1669390400
transform -1 0 49952 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _182_
timestamp 1669390400
transform -1 0 48496 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _183_
timestamp 1669390400
transform -1 0 46816 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _184_
timestamp 1669390400
transform 1 0 43568 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _185_
timestamp 1669390400
transform 1 0 43680 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _186_
timestamp 1669390400
transform 1 0 53872 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1669390400
transform -1 0 46928 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1669390400
transform -1 0 45024 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1669390400
transform 1 0 44352 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1669390400
transform -1 0 46144 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _191_
timestamp 1669390400
transform -1 0 46144 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1669390400
transform -1 0 45808 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1669390400
transform 1 0 45360 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _194_
timestamp 1669390400
transform 1 0 44240 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _195_
timestamp 1669390400
transform 1 0 43568 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _196_
timestamp 1669390400
transform 1 0 51744 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _197_
timestamp 1669390400
transform 1 0 44016 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _198_
timestamp 1669390400
transform -1 0 48944 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _199_
timestamp 1669390400
transform 1 0 41440 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 56560 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1669390400
transform -1 0 58240 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1669390400
transform 1 0 47040 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1669390400
transform -1 0 58240 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _204_ ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 39872 0 1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _205_
timestamp 1669390400
transform -1 0 58240 0 1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1669390400
transform 1 0 45360 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1669390400
transform -1 0 56560 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1669390400
transform -1 0 53872 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1669390400
transform 1 0 41440 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1669390400
transform -1 0 43008 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1669390400
transform -1 0 58240 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1669390400
transform -1 0 53200 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1669390400
transform 1 0 47376 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1669390400
transform 1 0 54992 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1669390400
transform -1 0 43568 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1669390400
transform -1 0 42672 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1669390400
transform 1 0 54992 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1669390400
transform 1 0 52640 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1669390400
transform -1 0 44688 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout22 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 55664 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout23 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54768 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout24 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 55440 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1
timestamp 1669390400
transform -1 0 56560 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 54768 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform 1 0 5600 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform 1 0 54320 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform 1 0 29120 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform -1 0 56560 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input7
timestamp 1669390400
transform 1 0 45808 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input8
timestamp 1669390400
transform -1 0 56560 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input9
timestamp 1669390400
transform -1 0 56560 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform 1 0 11200 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 56560 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output12 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3248 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output13
timestamp 1669390400
transform 1 0 54768 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output14
timestamp 1669390400
transform -1 0 3248 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output15
timestamp 1669390400
transform -1 0 50736 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output16
timestamp 1669390400
transform -1 0 56336 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output17
timestamp 1669390400
transform -1 0 3248 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18
timestamp 1669390400
transform -1 0 4368 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 56336 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform 1 0 56560 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform -1 0 12992 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_25 ~/sky130/gf180/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 57792 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_26
timestamp 1669390400
transform -1 0 22736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_27
timestamp 1669390400
transform -1 0 2128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_28
timestamp 1669390400
transform -1 0 2128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_29
timestamp 1669390400
transform -1 0 2128 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_30
timestamp 1669390400
transform -1 0 39536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_31
timestamp 1669390400
transform -1 0 5152 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_32
timestamp 1669390400
transform -1 0 37408 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_33
timestamp 1669390400
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_34
timestamp 1669390400
transform -1 0 2128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_35
timestamp 1669390400
transform 1 0 57792 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_36
timestamp 1669390400
transform -1 0 2128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_37
timestamp 1669390400
transform -1 0 16688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_38
timestamp 1669390400
transform -1 0 2800 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_39
timestamp 1669390400
transform 1 0 57792 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_40
timestamp 1669390400
transform -1 0 2128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_41
timestamp 1669390400
transform 1 0 55664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_42
timestamp 1669390400
transform -1 0 27440 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_43
timestamp 1669390400
transform 1 0 10752 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_44
timestamp 1669390400
transform -1 0 2128 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_45
timestamp 1669390400
transform -1 0 58240 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_46
timestamp 1669390400
transform -1 0 2128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_47
timestamp 1669390400
transform -1 0 2128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_48
timestamp 1669390400
transform -1 0 15344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_49
timestamp 1669390400
transform -1 0 58240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_50
timestamp 1669390400
transform -1 0 2800 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_51
timestamp 1669390400
transform 1 0 57792 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_52
timestamp 1669390400
transform -1 0 2128 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_53
timestamp 1669390400
transform -1 0 47600 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_54
timestamp 1669390400
transform -1 0 22736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_55
timestamp 1669390400
transform -1 0 2128 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_56
timestamp 1669390400
transform -1 0 28672 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_57
timestamp 1669390400
transform -1 0 3920 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_58
timestamp 1669390400
transform 1 0 57792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_59
timestamp 1669390400
transform -1 0 57008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_60
timestamp 1669390400
transform -1 0 38864 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_61
timestamp 1669390400
transform 1 0 47824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_62
timestamp 1669390400
transform -1 0 2800 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_63
timestamp 1669390400
transform -1 0 14672 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_64
timestamp 1669390400
transform -1 0 49840 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_65
timestamp 1669390400
transform -1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_66
timestamp 1669390400
transform 1 0 57792 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_67
timestamp 1669390400
transform -1 0 9968 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_68
timestamp 1669390400
transform 1 0 57792 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_69
timestamp 1669390400
transform -1 0 3472 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_70
timestamp 1669390400
transform -1 0 2128 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_71
timestamp 1669390400
transform 1 0 57792 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_72
timestamp 1669390400
transform 1 0 57792 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_73
timestamp 1669390400
transform -1 0 2128 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_74
timestamp 1669390400
transform -1 0 52080 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_75
timestamp 1669390400
transform 1 0 57120 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_76
timestamp 1669390400
transform -1 0 2128 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_77
timestamp 1669390400
transform 1 0 57792 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_78
timestamp 1669390400
transform -1 0 2128 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_79
timestamp 1669390400
transform -1 0 19376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_80
timestamp 1669390400
transform -1 0 2128 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_81
timestamp 1669390400
transform 1 0 57792 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_82
timestamp 1669390400
transform -1 0 14000 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_83
timestamp 1669390400
transform 1 0 57792 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_84
timestamp 1669390400
transform -1 0 2128 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_85
timestamp 1669390400
transform -1 0 32144 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_86
timestamp 1669390400
transform -1 0 3920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_87
timestamp 1669390400
transform -1 0 51408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_88
timestamp 1669390400
transform -1 0 2128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_89
timestamp 1669390400
transform -1 0 4592 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_90
timestamp 1669390400
transform -1 0 24752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_91
timestamp 1669390400
transform -1 0 42000 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_92
timestamp 1669390400
transform 1 0 57792 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_93
timestamp 1669390400
transform -1 0 14000 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_94
timestamp 1669390400
transform 1 0 57120 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_95
timestamp 1669390400
transform -1 0 2128 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_96
timestamp 1669390400
transform -1 0 2128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_97
timestamp 1669390400
transform -1 0 38080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_98
timestamp 1669390400
transform -1 0 21728 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_99
timestamp 1669390400
transform -1 0 2128 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_100
timestamp 1669390400
transform -1 0 30128 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_101
timestamp 1669390400
transform -1 0 34160 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_102
timestamp 1669390400
transform 1 0 57792 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_103
timestamp 1669390400
transform -1 0 2128 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_104
timestamp 1669390400
transform -1 0 46928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_105
timestamp 1669390400
transform 1 0 57792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_106
timestamp 1669390400
transform -1 0 13888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_107
timestamp 1669390400
transform -1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_108
timestamp 1669390400
transform -1 0 2128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_109
timestamp 1669390400
transform 1 0 57792 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_110
timestamp 1669390400
transform -1 0 37408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_111
timestamp 1669390400
transform -1 0 41328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_112
timestamp 1669390400
transform -1 0 39536 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_113
timestamp 1669390400
transform 1 0 57792 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_114
timestamp 1669390400
transform -1 0 2128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_115
timestamp 1669390400
transform 1 0 57792 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_116
timestamp 1669390400
transform -1 0 49168 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_117
timestamp 1669390400
transform 1 0 57792 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_118
timestamp 1669390400
transform -1 0 48272 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_119
timestamp 1669390400
transform -1 0 2128 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_120
timestamp 1669390400
transform -1 0 2128 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_121
timestamp 1669390400
transform -1 0 40208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_122
timestamp 1669390400
transform -1 0 2800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_123
timestamp 1669390400
transform -1 0 2128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_124
timestamp 1669390400
transform -1 0 2128 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_125
timestamp 1669390400
transform -1 0 19376 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_126
timestamp 1669390400
transform -1 0 2128 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_127
timestamp 1669390400
transform -1 0 12656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_128
timestamp 1669390400
transform -1 0 4592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_129
timestamp 1669390400
transform -1 0 33488 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_130
timestamp 1669390400
transform -1 0 20048 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_131
timestamp 1669390400
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_132
timestamp 1669390400
transform -1 0 44240 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_133
timestamp 1669390400
transform -1 0 2800 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  top_wrapper_134
timestamp 1669390400
transform 1 0 57792 0 1 45472
box -86 -86 534 870
<< labels >>
flabel metal3 s 59200 36904 59800 37128 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 59200 48328 59800 48552 0 FreeSans 896 0 0 0 io_in[1]
port 1 nsew signal input
flabel metal2 s 5320 59200 5544 59800 0 FreeSans 896 90 0 0 io_in[2]
port 2 nsew signal input
flabel metal2 s 58408 59200 58632 59800 0 FreeSans 896 90 0 0 io_in[3]
port 3 nsew signal input
flabel metal2 s 28168 200 28392 800 0 FreeSans 896 90 0 0 io_in[4]
port 4 nsew signal input
flabel metal3 s 59200 22792 59800 23016 0 FreeSans 896 0 0 0 io_in[5]
port 5 nsew signal input
flabel metal2 s 45640 59200 45864 59800 0 FreeSans 896 90 0 0 io_in[6]
port 6 nsew signal input
flabel metal2 s 59080 59200 59304 59800 0 FreeSans 896 90 0 0 io_in[7]
port 7 nsew signal input
flabel metal3 s 59200 19432 59800 19656 0 FreeSans 896 0 0 0 io_in[8]
port 8 nsew signal input
flabel metal2 s 11368 200 11592 800 0 FreeSans 896 90 0 0 io_in[9]
port 9 nsew signal input
flabel metal3 s 59200 52360 59800 52584 0 FreeSans 896 0 0 0 io_oeb[0]
port 10 nsew signal tristate
flabel metal2 s 22120 59200 22344 59800 0 FreeSans 896 90 0 0 io_oeb[1]
port 11 nsew signal tristate
flabel metal3 s 200 1960 800 2184 0 FreeSans 896 0 0 0 io_oeb[2]
port 12 nsew signal tristate
flabel metal3 s 200 14056 800 14280 0 FreeSans 896 0 0 0 io_oeb[3]
port 13 nsew signal tristate
flabel metal3 s 200 39592 800 39816 0 FreeSans 896 0 0 0 io_oeb[4]
port 14 nsew signal tristate
flabel metal2 s 38920 200 39144 800 0 FreeSans 896 90 0 0 io_oeb[5]
port 15 nsew signal tristate
flabel metal2 s 4648 59200 4872 59800 0 FreeSans 896 90 0 0 io_oeb[6]
port 16 nsew signal tristate
flabel metal2 s 36232 59200 36456 59800 0 FreeSans 896 90 0 0 io_oeb[7]
port 17 nsew signal tristate
flabel metal2 s 34888 200 35112 800 0 FreeSans 896 90 0 0 io_oeb[8]
port 18 nsew signal tristate
flabel metal3 s 200 12712 800 12936 0 FreeSans 896 0 0 0 io_oeb[9]
port 19 nsew signal tristate
flabel metal3 s 200 53032 800 53256 0 FreeSans 896 0 0 0 io_out[0]
port 20 nsew signal tristate
flabel metal3 s 59200 40936 59800 41160 0 FreeSans 896 0 0 0 io_out[1]
port 21 nsew signal tristate
flabel metal3 s 200 54376 800 54600 0 FreeSans 896 0 0 0 io_out[2]
port 22 nsew signal tristate
flabel metal2 s 49000 200 49224 800 0 FreeSans 896 90 0 0 io_out[3]
port 23 nsew signal tristate
flabel metal3 s 59200 49672 59800 49896 0 FreeSans 896 0 0 0 io_out[4]
port 24 nsew signal tristate
flabel metal3 s 200 24808 800 25032 0 FreeSans 896 0 0 0 io_out[5]
port 25 nsew signal tristate
flabel metal2 s 2632 59200 2856 59800 0 FreeSans 896 90 0 0 io_out[6]
port 26 nsew signal tristate
flabel metal3 s 59200 34888 59800 35112 0 FreeSans 896 0 0 0 io_out[7]
port 27 nsew signal tristate
flabel metal2 s 56392 59200 56616 59800 0 FreeSans 896 90 0 0 io_out[8]
port 28 nsew signal tristate
flabel metal2 s 12040 59200 12264 59800 0 FreeSans 896 90 0 0 io_out[9]
port 29 nsew signal tristate
flabel metal3 s 59200 26824 59800 27048 0 FreeSans 896 0 0 0 la_data_in[0]
port 30 nsew signal input
flabel metal2 s 20776 200 21000 800 0 FreeSans 896 90 0 0 la_data_in[10]
port 31 nsew signal input
flabel metal3 s 59200 4648 59800 4872 0 FreeSans 896 0 0 0 la_data_in[11]
port 32 nsew signal input
flabel metal3 s 59200 22120 59800 22344 0 FreeSans 896 0 0 0 la_data_in[12]
port 33 nsew signal input
flabel metal2 s 57064 59200 57288 59800 0 FreeSans 896 90 0 0 la_data_in[13]
port 34 nsew signal input
flabel metal2 s 29512 200 29736 800 0 FreeSans 896 90 0 0 la_data_in[14]
port 35 nsew signal input
flabel metal3 s 59200 24808 59800 25032 0 FreeSans 896 0 0 0 la_data_in[15]
port 36 nsew signal input
flabel metal2 s 616 59200 840 59800 0 FreeSans 896 90 0 0 la_data_in[16]
port 37 nsew signal input
flabel metal3 s 200 59080 800 59304 0 FreeSans 896 0 0 0 la_data_in[17]
port 38 nsew signal input
flabel metal2 s 17416 200 17640 800 0 FreeSans 896 90 0 0 la_data_in[18]
port 39 nsew signal input
flabel metal2 s 44968 200 45192 800 0 FreeSans 896 90 0 0 la_data_in[19]
port 40 nsew signal input
flabel metal2 s 44968 59200 45192 59800 0 FreeSans 896 90 0 0 la_data_in[1]
port 41 nsew signal input
flabel metal2 s 22792 59200 23016 59800 0 FreeSans 896 90 0 0 la_data_in[20]
port 42 nsew signal input
flabel metal3 s 59200 26152 59800 26376 0 FreeSans 896 0 0 0 la_data_in[21]
port 43 nsew signal input
flabel metal3 s 200 27496 800 27720 0 FreeSans 896 0 0 0 la_data_in[22]
port 44 nsew signal input
flabel metal2 s 10024 59200 10248 59800 0 FreeSans 896 90 0 0 la_data_in[23]
port 45 nsew signal input
flabel metal2 s 23464 200 23688 800 0 FreeSans 896 90 0 0 la_data_in[24]
port 46 nsew signal input
flabel metal2 s 28840 59200 29064 59800 0 FreeSans 896 90 0 0 la_data_in[25]
port 47 nsew signal input
flabel metal3 s 59200 41608 59800 41832 0 FreeSans 896 0 0 0 la_data_in[26]
port 48 nsew signal input
flabel metal2 s 53032 59200 53256 59800 0 FreeSans 896 90 0 0 la_data_in[27]
port 49 nsew signal input
flabel metal3 s 200 23464 800 23688 0 FreeSans 896 0 0 0 la_data_in[28]
port 50 nsew signal input
flabel metal3 s 59200 6664 59800 6888 0 FreeSans 896 0 0 0 la_data_in[29]
port 51 nsew signal input
flabel metal3 s 200 55720 800 55944 0 FreeSans 896 0 0 0 la_data_in[2]
port 52 nsew signal input
flabel metal3 s 59200 56392 59800 56616 0 FreeSans 896 0 0 0 la_data_in[30]
port 53 nsew signal input
flabel metal3 s 59200 37576 59800 37800 0 FreeSans 896 0 0 0 la_data_in[31]
port 54 nsew signal input
flabel metal3 s 200 41608 800 41832 0 FreeSans 896 0 0 0 la_data_in[32]
port 55 nsew signal input
flabel metal2 s 55048 200 55272 800 0 FreeSans 896 90 0 0 la_data_in[33]
port 56 nsew signal input
flabel metal3 s 59200 9352 59800 9576 0 FreeSans 896 0 0 0 la_data_in[34]
port 57 nsew signal input
flabel metal2 s 49672 59200 49896 59800 0 FreeSans 896 90 0 0 la_data_in[35]
port 58 nsew signal input
flabel metal2 s 7336 59200 7560 59800 0 FreeSans 896 90 0 0 la_data_in[36]
port 59 nsew signal input
flabel metal2 s 52360 59200 52584 59800 0 FreeSans 896 90 0 0 la_data_in[37]
port 60 nsew signal input
flabel metal3 s 200 37576 800 37800 0 FreeSans 896 0 0 0 la_data_in[38]
port 61 nsew signal input
flabel metal2 s 14728 59200 14952 59800 0 FreeSans 896 90 0 0 la_data_in[39]
port 62 nsew signal input
flabel metal3 s 200 2632 800 2856 0 FreeSans 896 0 0 0 la_data_in[3]
port 63 nsew signal input
flabel metal2 s 26152 59200 26376 59800 0 FreeSans 896 90 0 0 la_data_in[40]
port 64 nsew signal input
flabel metal2 s 15400 200 15624 800 0 FreeSans 896 90 0 0 la_data_in[41]
port 65 nsew signal input
flabel metal3 s 59200 10024 59800 10248 0 FreeSans 896 0 0 0 la_data_in[42]
port 66 nsew signal input
flabel metal2 s 54376 59200 54600 59800 0 FreeSans 896 90 0 0 la_data_in[43]
port 67 nsew signal input
flabel metal2 s 33544 200 33768 800 0 FreeSans 896 90 0 0 la_data_in[44]
port 68 nsew signal input
flabel metal3 s 59200 38248 59800 38472 0 FreeSans 896 0 0 0 la_data_in[45]
port 69 nsew signal input
flabel metal3 s 200 6664 800 6888 0 FreeSans 896 0 0 0 la_data_in[46]
port 70 nsew signal input
flabel metal3 s 59200 5992 59800 6216 0 FreeSans 896 0 0 0 la_data_in[47]
port 71 nsew signal input
flabel metal2 s 27496 200 27720 800 0 FreeSans 896 90 0 0 la_data_in[48]
port 72 nsew signal input
flabel metal3 s 200 12040 800 12264 0 FreeSans 896 0 0 0 la_data_in[49]
port 73 nsew signal input
flabel metal3 s 200 42280 800 42504 0 FreeSans 896 0 0 0 la_data_in[4]
port 74 nsew signal input
flabel metal3 s 200 3304 800 3528 0 FreeSans 896 0 0 0 la_data_in[50]
port 75 nsew signal input
flabel metal3 s 200 32200 800 32424 0 FreeSans 896 0 0 0 la_data_in[51]
port 76 nsew signal input
flabel metal2 s 17416 59200 17640 59800 0 FreeSans 896 90 0 0 la_data_in[52]
port 77 nsew signal input
flabel metal3 s 59200 2632 59800 2856 0 FreeSans 896 0 0 0 la_data_in[53]
port 78 nsew signal input
flabel metal3 s 59200 14056 59800 14280 0 FreeSans 896 0 0 0 la_data_in[54]
port 79 nsew signal input
flabel metal3 s 200 20104 800 20328 0 FreeSans 896 0 0 0 la_data_in[55]
port 80 nsew signal input
flabel metal2 s 24808 200 25032 800 0 FreeSans 896 90 0 0 la_data_in[56]
port 81 nsew signal input
flabel metal2 s 38248 200 38472 800 0 FreeSans 896 90 0 0 la_data_in[57]
port 82 nsew signal input
flabel metal2 s 21448 59200 21672 59800 0 FreeSans 896 90 0 0 la_data_in[58]
port 83 nsew signal input
flabel metal3 s 59200 55048 59800 55272 0 FreeSans 896 0 0 0 la_data_in[59]
port 84 nsew signal input
flabel metal2 s 24136 59200 24360 59800 0 FreeSans 896 90 0 0 la_data_in[5]
port 85 nsew signal input
flabel metal2 s 56392 200 56616 800 0 FreeSans 896 90 0 0 la_data_in[60]
port 86 nsew signal input
flabel metal2 s 19432 200 19656 800 0 FreeSans 896 90 0 0 la_data_in[61]
port 87 nsew signal input
flabel metal3 s 200 33544 800 33768 0 FreeSans 896 0 0 0 la_data_in[62]
port 88 nsew signal input
flabel metal3 s 59200 11368 59800 11592 0 FreeSans 896 0 0 0 la_data_in[63]
port 89 nsew signal input
flabel metal2 s 7336 200 7560 800 0 FreeSans 896 90 0 0 la_data_in[6]
port 90 nsew signal input
flabel metal2 s 6664 59200 6888 59800 0 FreeSans 896 90 0 0 la_data_in[7]
port 91 nsew signal input
flabel metal2 s 15400 59200 15624 59800 0 FreeSans 896 90 0 0 la_data_in[8]
port 92 nsew signal input
flabel metal3 s 200 7336 800 7560 0 FreeSans 896 0 0 0 la_data_in[9]
port 93 nsew signal input
flabel metal3 s 59200 -56 59800 168 0 FreeSans 896 0 0 0 la_data_out[0]
port 94 nsew signal tristate
flabel metal2 s 57736 59200 57960 59800 0 FreeSans 896 90 0 0 la_data_out[10]
port 95 nsew signal tristate
flabel metal3 s 200 26824 800 27048 0 FreeSans 896 0 0 0 la_data_out[11]
port 96 nsew signal tristate
flabel metal3 s 200 21448 800 21672 0 FreeSans 896 0 0 0 la_data_out[12]
port 97 nsew signal tristate
flabel metal2 s 14728 200 14952 800 0 FreeSans 896 90 0 0 la_data_out[13]
port 98 nsew signal tristate
flabel metal2 s 57736 200 57960 800 0 FreeSans 896 90 0 0 la_data_out[14]
port 99 nsew signal tristate
flabel metal3 s 200 45640 800 45864 0 FreeSans 896 0 0 0 la_data_out[15]
port 100 nsew signal tristate
flabel metal3 s 59200 3304 59800 3528 0 FreeSans 896 0 0 0 la_data_out[16]
port 101 nsew signal tristate
flabel metal3 s 200 44296 800 44520 0 FreeSans 896 0 0 0 la_data_out[17]
port 102 nsew signal tristate
flabel metal2 s 46984 200 47208 800 0 FreeSans 896 90 0 0 la_data_out[18]
port 103 nsew signal tristate
flabel metal2 s 22120 200 22344 800 0 FreeSans 896 90 0 0 la_data_out[19]
port 104 nsew signal tristate
flabel metal3 s 200 28168 800 28392 0 FreeSans 896 0 0 0 la_data_out[1]
port 105 nsew signal tristate
flabel metal3 s 200 34888 800 35112 0 FreeSans 896 0 0 0 la_data_out[20]
port 106 nsew signal tristate
flabel metal2 s 28168 59200 28392 59800 0 FreeSans 896 90 0 0 la_data_out[21]
port 107 nsew signal tristate
flabel metal2 s 3304 59200 3528 59800 0 FreeSans 896 90 0 0 la_data_out[22]
port 108 nsew signal tristate
flabel metal3 s 59200 28168 59800 28392 0 FreeSans 896 0 0 0 la_data_out[23]
port 109 nsew signal tristate
flabel metal2 s 55720 200 55944 800 0 FreeSans 896 90 0 0 la_data_out[24]
port 110 nsew signal tristate
flabel metal2 s 38248 59200 38472 59800 0 FreeSans 896 90 0 0 la_data_out[25]
port 111 nsew signal tristate
flabel metal2 s 48328 200 48552 800 0 FreeSans 896 90 0 0 la_data_out[26]
port 112 nsew signal tristate
flabel metal2 s 1288 59200 1512 59800 0 FreeSans 896 90 0 0 la_data_out[27]
port 113 nsew signal tristate
flabel metal2 s 14056 59200 14280 59800 0 FreeSans 896 90 0 0 la_data_out[28]
port 114 nsew signal tristate
flabel metal2 s 49000 59200 49224 59800 0 FreeSans 896 90 0 0 la_data_out[29]
port 115 nsew signal tristate
flabel metal2 s 16072 200 16296 800 0 FreeSans 896 90 0 0 la_data_out[2]
port 116 nsew signal tristate
flabel metal2 s 16072 59200 16296 59800 0 FreeSans 896 90 0 0 la_data_out[30]
port 117 nsew signal tristate
flabel metal3 s 59200 30184 59800 30408 0 FreeSans 896 0 0 0 la_data_out[31]
port 118 nsew signal tristate
flabel metal2 s 9352 59200 9576 59800 0 FreeSans 896 90 0 0 la_data_out[32]
port 119 nsew signal tristate
flabel metal3 s 59200 40264 59800 40488 0 FreeSans 896 0 0 0 la_data_out[33]
port 120 nsew signal tristate
flabel metal3 s 200 58408 800 58632 0 FreeSans 896 0 0 0 la_data_out[34]
port 121 nsew signal tristate
flabel metal3 s 200 46984 800 47208 0 FreeSans 896 0 0 0 la_data_out[35]
port 122 nsew signal tristate
flabel metal3 s 59200 46312 59800 46536 0 FreeSans 896 0 0 0 la_data_out[36]
port 123 nsew signal tristate
flabel metal3 s 59200 51016 59800 51240 0 FreeSans 896 0 0 0 la_data_out[37]
port 124 nsew signal tristate
flabel metal3 s 200 19432 800 19656 0 FreeSans 896 0 0 0 la_data_out[38]
port 125 nsew signal tristate
flabel metal2 s 51016 200 51240 800 0 FreeSans 896 90 0 0 la_data_out[39]
port 126 nsew signal tristate
flabel metal3 s 200 30856 800 31080 0 FreeSans 896 0 0 0 la_data_out[3]
port 127 nsew signal tristate
flabel metal3 s 59200 58408 59800 58632 0 FreeSans 896 0 0 0 la_data_out[40]
port 128 nsew signal tristate
flabel metal3 s 200 51016 800 51240 0 FreeSans 896 0 0 0 la_data_out[41]
port 129 nsew signal tristate
flabel metal3 s 59200 24136 59800 24360 0 FreeSans 896 0 0 0 la_data_out[42]
port 130 nsew signal tristate
flabel metal3 s 200 53704 800 53928 0 FreeSans 896 0 0 0 la_data_out[43]
port 131 nsew signal tristate
flabel metal2 s 18760 200 18984 800 0 FreeSans 896 90 0 0 la_data_out[44]
port 132 nsew signal tristate
flabel metal3 s 200 4648 800 4872 0 FreeSans 896 0 0 0 la_data_out[45]
port 133 nsew signal tristate
flabel metal3 s 59200 38920 59800 39144 0 FreeSans 896 0 0 0 la_data_out[46]
port 134 nsew signal tristate
flabel metal2 s 13384 59200 13608 59800 0 FreeSans 896 90 0 0 la_data_out[47]
port 135 nsew signal tristate
flabel metal2 s 59752 59200 59976 59800 0 FreeSans 896 90 0 0 la_data_out[48]
port 136 nsew signal tristate
flabel metal3 s 200 18088 800 18312 0 FreeSans 896 0 0 0 la_data_out[49]
port 137 nsew signal tristate
flabel metal3 s 59200 10696 59800 10920 0 FreeSans 896 0 0 0 la_data_out[4]
port 138 nsew signal tristate
flabel metal2 s 31528 59200 31752 59800 0 FreeSans 896 90 0 0 la_data_out[50]
port 139 nsew signal tristate
flabel metal2 s 3304 200 3528 800 0 FreeSans 896 90 0 0 la_data_out[51]
port 140 nsew signal tristate
flabel metal2 s 50344 200 50568 800 0 FreeSans 896 90 0 0 la_data_out[52]
port 141 nsew signal tristate
flabel metal3 s 200 44968 800 45192 0 FreeSans 896 0 0 0 la_data_out[53]
port 142 nsew signal tristate
flabel metal3 s 200 57064 800 57288 0 FreeSans 896 0 0 0 la_data_out[54]
port 143 nsew signal tristate
flabel metal2 s 24136 200 24360 800 0 FreeSans 896 90 0 0 la_data_out[55]
port 144 nsew signal tristate
flabel metal2 s 40936 59200 41160 59800 0 FreeSans 896 90 0 0 la_data_out[56]
port 145 nsew signal tristate
flabel metal3 s 59200 47656 59800 47880 0 FreeSans 896 0 0 0 la_data_out[57]
port 146 nsew signal tristate
flabel metal2 s 12712 59200 12936 59800 0 FreeSans 896 90 0 0 la_data_out[58]
port 147 nsew signal tristate
flabel metal3 s 59200 30856 59800 31080 0 FreeSans 896 0 0 0 la_data_out[59]
port 148 nsew signal tristate
flabel metal3 s 200 38920 800 39144 0 FreeSans 896 0 0 0 la_data_out[5]
port 149 nsew signal tristate
flabel metal3 s 200 10024 800 10248 0 FreeSans 896 0 0 0 la_data_out[60]
port 150 nsew signal tristate
flabel metal3 s 200 9352 800 9576 0 FreeSans 896 0 0 0 la_data_out[61]
port 151 nsew signal tristate
flabel metal2 s 36904 59200 37128 59800 0 FreeSans 896 90 0 0 la_data_out[62]
port 152 nsew signal tristate
flabel metal2 s 20776 59200 21000 59800 0 FreeSans 896 90 0 0 la_data_out[63]
port 153 nsew signal tristate
flabel metal3 s 59200 1960 59800 2184 0 FreeSans 896 0 0 0 la_data_out[6]
port 154 nsew signal tristate
flabel metal2 s 26824 59200 27048 59800 0 FreeSans 896 90 0 0 la_data_out[7]
port 155 nsew signal tristate
flabel metal2 s 11368 59200 11592 59800 0 FreeSans 896 90 0 0 la_data_out[8]
port 156 nsew signal tristate
flabel metal3 s 200 52360 800 52584 0 FreeSans 896 0 0 0 la_data_out[9]
port 157 nsew signal tristate
flabel metal3 s 59200 7336 59800 7560 0 FreeSans 896 0 0 0 la_oenb[0]
port 158 nsew signal input
flabel metal3 s 200 30184 800 30408 0 FreeSans 896 0 0 0 la_oenb[10]
port 159 nsew signal input
flabel metal3 s 59200 17416 59800 17640 0 FreeSans 896 0 0 0 la_oenb[11]
port 160 nsew signal input
flabel metal2 s 37576 200 37800 800 0 FreeSans 896 90 0 0 la_oenb[12]
port 161 nsew signal input
flabel metal2 s 34888 59200 35112 59800 0 FreeSans 896 90 0 0 la_oenb[13]
port 162 nsew signal input
flabel metal2 s 36904 200 37128 800 0 FreeSans 896 90 0 0 la_oenb[14]
port 163 nsew signal input
flabel metal3 s 200 1288 800 1512 0 FreeSans 896 0 0 0 la_oenb[15]
port 164 nsew signal input
flabel metal2 s 6664 200 6888 800 0 FreeSans 896 90 0 0 la_oenb[16]
port 165 nsew signal input
flabel metal2 s 10696 200 10920 800 0 FreeSans 896 90 0 0 la_oenb[17]
port 166 nsew signal input
flabel metal2 s 44296 59200 44520 59800 0 FreeSans 896 90 0 0 la_oenb[18]
port 167 nsew signal input
flabel metal2 s 42280 59200 42504 59800 0 FreeSans 896 90 0 0 la_oenb[19]
port 168 nsew signal input
flabel metal3 s 200 11368 800 11592 0 FreeSans 896 0 0 0 la_oenb[1]
port 169 nsew signal input
flabel metal3 s 59200 44968 59800 45192 0 FreeSans 896 0 0 0 la_oenb[20]
port 170 nsew signal input
flabel metal3 s 200 5320 800 5544 0 FreeSans 896 0 0 0 la_oenb[21]
port 171 nsew signal input
flabel metal3 s 200 36904 800 37128 0 FreeSans 896 0 0 0 la_oenb[22]
port 172 nsew signal input
flabel metal2 s 14056 200 14280 800 0 FreeSans 896 90 0 0 la_oenb[23]
port 173 nsew signal input
flabel metal2 s 23464 59200 23688 59800 0 FreeSans 896 90 0 0 la_oenb[24]
port 174 nsew signal input
flabel metal2 s 3976 59200 4200 59800 0 FreeSans 896 90 0 0 la_oenb[25]
port 175 nsew signal input
flabel metal3 s 200 10696 800 10920 0 FreeSans 896 0 0 0 la_oenb[26]
port 176 nsew signal input
flabel metal3 s 200 18760 800 18984 0 FreeSans 896 0 0 0 la_oenb[27]
port 177 nsew signal input
flabel metal3 s 59200 18088 59800 18312 0 FreeSans 896 0 0 0 la_oenb[28]
port 178 nsew signal input
flabel metal3 s 59200 39592 59800 39816 0 FreeSans 896 0 0 0 la_oenb[29]
port 179 nsew signal input
flabel metal3 s 59200 43624 59800 43848 0 FreeSans 896 0 0 0 la_oenb[2]
port 180 nsew signal input
flabel metal3 s 59200 35560 59800 35784 0 FreeSans 896 0 0 0 la_oenb[30]
port 181 nsew signal input
flabel metal2 s 47656 59200 47880 59800 0 FreeSans 896 90 0 0 la_oenb[31]
port 182 nsew signal input
flabel metal3 s 59200 33544 59800 33768 0 FreeSans 896 0 0 0 la_oenb[32]
port 183 nsew signal input
flabel metal2 s 26152 200 26376 800 0 FreeSans 896 90 0 0 la_oenb[33]
port 184 nsew signal input
flabel metal3 s 59200 49000 59800 49224 0 FreeSans 896 0 0 0 la_oenb[34]
port 185 nsew signal input
flabel metal3 s 200 26152 800 26376 0 FreeSans 896 0 0 0 la_oenb[35]
port 186 nsew signal input
flabel metal2 s 616 200 840 800 0 FreeSans 896 90 0 0 la_oenb[36]
port 187 nsew signal input
flabel metal2 s 35560 59200 35784 59800 0 FreeSans 896 90 0 0 la_oenb[37]
port 188 nsew signal input
flabel metal2 s 26824 200 27048 800 0 FreeSans 896 90 0 0 la_oenb[38]
port 189 nsew signal input
flabel metal2 s 54376 200 54600 800 0 FreeSans 896 90 0 0 la_oenb[39]
port 190 nsew signal input
flabel metal3 s 200 50344 800 50568 0 FreeSans 896 0 0 0 la_oenb[3]
port 191 nsew signal input
flabel metal2 s 58408 200 58632 800 0 FreeSans 896 90 0 0 la_oenb[40]
port 192 nsew signal input
flabel metal2 s 41608 59200 41832 59800 0 FreeSans 896 90 0 0 la_oenb[41]
port 193 nsew signal input
flabel metal3 s 200 47656 800 47880 0 FreeSans 896 0 0 0 la_oenb[42]
port 194 nsew signal input
flabel metal2 s 10024 200 10248 800 0 FreeSans 896 90 0 0 la_oenb[43]
port 195 nsew signal input
flabel metal3 s 200 8680 800 8904 0 FreeSans 896 0 0 0 la_oenb[44]
port 196 nsew signal input
flabel metal3 s 59200 54376 59800 54600 0 FreeSans 896 0 0 0 la_oenb[45]
port 197 nsew signal input
flabel metal2 s 41608 200 41832 800 0 FreeSans 896 90 0 0 la_oenb[46]
port 198 nsew signal input
flabel metal2 s 20104 200 20328 800 0 FreeSans 896 90 0 0 la_oenb[47]
port 199 nsew signal input
flabel metal3 s 200 32872 800 33096 0 FreeSans 896 0 0 0 la_oenb[48]
port 200 nsew signal input
flabel metal3 s 59200 18760 59800 18984 0 FreeSans 896 0 0 0 la_oenb[49]
port 201 nsew signal input
flabel metal2 s 8680 59200 8904 59800 0 FreeSans 896 90 0 0 la_oenb[4]
port 202 nsew signal input
flabel metal2 s 40936 200 41160 800 0 FreeSans 896 90 0 0 la_oenb[50]
port 203 nsew signal input
flabel metal2 s 37576 59200 37800 59800 0 FreeSans 896 90 0 0 la_oenb[51]
port 204 nsew signal input
flabel metal2 s 53032 200 53256 800 0 FreeSans 896 90 0 0 la_oenb[52]
port 205 nsew signal input
flabel metal3 s 200 46312 800 46536 0 FreeSans 896 0 0 0 la_oenb[53]
port 206 nsew signal input
flabel metal3 s 200 48328 800 48552 0 FreeSans 896 0 0 0 la_oenb[54]
port 207 nsew signal input
flabel metal3 s 59200 20776 59800 21000 0 FreeSans 896 0 0 0 la_oenb[55]
port 208 nsew signal input
flabel metal2 s 40264 200 40488 800 0 FreeSans 896 90 0 0 la_oenb[56]
port 209 nsew signal input
flabel metal3 s 59200 53704 59800 53928 0 FreeSans 896 0 0 0 la_oenb[57]
port 210 nsew signal input
flabel metal2 s 59080 200 59304 800 0 FreeSans 896 90 0 0 la_oenb[58]
port 211 nsew signal input
flabel metal2 s 50344 59200 50568 59800 0 FreeSans 896 90 0 0 la_oenb[59]
port 212 nsew signal input
flabel metal2 s 49672 200 49896 800 0 FreeSans 896 90 0 0 la_oenb[5]
port 213 nsew signal input
flabel metal2 s 30856 59200 31080 59800 0 FreeSans 896 90 0 0 la_oenb[60]
port 214 nsew signal input
flabel metal2 s 5992 200 6216 800 0 FreeSans 896 90 0 0 la_oenb[61]
port 215 nsew signal input
flabel metal3 s 59200 21448 59800 21672 0 FreeSans 896 0 0 0 la_oenb[62]
port 216 nsew signal input
flabel metal2 s 1960 59200 2184 59800 0 FreeSans 896 90 0 0 la_oenb[63]
port 217 nsew signal input
flabel metal3 s 200 616 800 840 0 FreeSans 896 0 0 0 la_oenb[6]
port 218 nsew signal input
flabel metal2 s 13384 200 13608 800 0 FreeSans 896 90 0 0 la_oenb[7]
port 219 nsew signal input
flabel metal2 s 52360 200 52584 800 0 FreeSans 896 90 0 0 la_oenb[8]
port 220 nsew signal input
flabel metal2 s 32200 59200 32424 59800 0 FreeSans 896 90 0 0 la_oenb[9]
port 221 nsew signal input
flabel metal3 s 59200 57064 59800 57288 0 FreeSans 896 0 0 0 user_clock2
port 222 nsew signal input
flabel metal3 s 200 40264 800 40488 0 FreeSans 896 0 0 0 user_irq[0]
port 223 nsew signal tristate
flabel metal2 s 29512 59200 29736 59800 0 FreeSans 896 90 0 0 user_irq[1]
port 224 nsew signal tristate
flabel metal2 s 33544 59200 33768 59800 0 FreeSans 896 90 0 0 user_irq[2]
port 225 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 226 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 226 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 227 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 227 nsew ground bidirectional
flabel metal3 s 59200 3976 59800 4200 0 FreeSans 896 0 0 0 wb_clk_i
port 228 nsew signal input
flabel metal2 s 24808 59200 25032 59800 0 FreeSans 896 90 0 0 wb_rst_i
port 229 nsew signal input
flabel metal3 s 59200 13384 59800 13608 0 FreeSans 896 0 0 0 wbs_ack_o
port 230 nsew signal tristate
flabel metal3 s 200 29512 800 29736 0 FreeSans 896 0 0 0 wbs_adr_i[0]
port 231 nsew signal input
flabel metal2 s 39592 59200 39816 59800 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 232 nsew signal input
flabel metal2 s 18088 59200 18312 59800 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 233 nsew signal input
flabel metal2 s 4648 200 4872 800 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 234 nsew signal input
flabel metal2 s 30856 200 31080 800 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 235 nsew signal input
flabel metal3 s 59200 36232 59800 36456 0 FreeSans 896 0 0 0 wbs_adr_i[14]
port 236 nsew signal input
flabel metal3 s 200 35560 800 35784 0 FreeSans 896 0 0 0 wbs_adr_i[15]
port 237 nsew signal input
flabel metal2 s 35560 200 35784 800 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 238 nsew signal input
flabel metal3 s 200 49000 800 49224 0 FreeSans 896 0 0 0 wbs_adr_i[17]
port 239 nsew signal input
flabel metal3 s 59200 12712 59800 12936 0 FreeSans 896 0 0 0 wbs_adr_i[18]
port 240 nsew signal input
flabel metal2 s 53704 200 53928 800 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 241 nsew signal input
flabel metal3 s 200 24136 800 24360 0 FreeSans 896 0 0 0 wbs_adr_i[1]
port 242 nsew signal input
flabel metal3 s 59200 55720 59800 55944 0 FreeSans 896 0 0 0 wbs_adr_i[20]
port 243 nsew signal input
flabel metal2 s 31528 200 31752 800 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 244 nsew signal input
flabel metal2 s 45640 200 45864 800 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 245 nsew signal input
flabel metal3 s 59200 8680 59800 8904 0 FreeSans 896 0 0 0 wbs_adr_i[23]
port 246 nsew signal input
flabel metal3 s 200 17416 800 17640 0 FreeSans 896 0 0 0 wbs_adr_i[24]
port 247 nsew signal input
flabel metal2 s 30184 200 30408 800 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 248 nsew signal input
flabel metal2 s 5320 200 5544 800 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 249 nsew signal input
flabel metal2 s 30184 59200 30408 59800 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 250 nsew signal input
flabel metal3 s 59200 28840 59800 29064 0 FreeSans 896 0 0 0 wbs_adr_i[28]
port 251 nsew signal input
flabel metal3 s 200 28840 800 29064 0 FreeSans 896 0 0 0 wbs_adr_i[29]
port 252 nsew signal input
flabel metal2 s 21448 200 21672 800 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 253 nsew signal input
flabel metal2 s 55720 59200 55944 59800 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 254 nsew signal input
flabel metal3 s 59200 20104 59800 20328 0 FreeSans 896 0 0 0 wbs_adr_i[31]
port 255 nsew signal input
flabel metal2 s 44296 200 44520 800 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 256 nsew signal input
flabel metal2 s 53704 59200 53928 59800 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 257 nsew signal input
flabel metal2 s 42280 200 42504 800 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 258 nsew signal input
flabel metal3 s 200 36232 800 36456 0 FreeSans 896 0 0 0 wbs_adr_i[6]
port 259 nsew signal input
flabel metal2 s 2632 200 2856 800 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 260 nsew signal input
flabel metal2 s 57064 200 57288 800 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 261 nsew signal input
flabel metal3 s 59200 12040 59800 12264 0 FreeSans 896 0 0 0 wbs_adr_i[9]
port 262 nsew signal input
flabel metal2 s 27496 59200 27720 59800 0 FreeSans 896 90 0 0 wbs_cyc_i
port 263 nsew signal input
flabel metal3 s 59200 46984 59800 47208 0 FreeSans 896 0 0 0 wbs_dat_i[0]
port 264 nsew signal input
flabel metal3 s 200 3976 800 4200 0 FreeSans 896 0 0 0 wbs_dat_i[10]
port 265 nsew signal input
flabel metal3 s 200 59752 800 59976 0 FreeSans 896 0 0 0 wbs_dat_i[11]
port 266 nsew signal input
flabel metal3 s 200 57736 800 57960 0 FreeSans 896 0 0 0 wbs_dat_i[12]
port 267 nsew signal input
flabel metal2 s 1960 200 2184 800 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 268 nsew signal input
flabel metal3 s 200 15400 800 15624 0 FreeSans 896 0 0 0 wbs_dat_i[14]
port 269 nsew signal input
flabel metal3 s 59200 27496 59800 27720 0 FreeSans 896 0 0 0 wbs_dat_i[15]
port 270 nsew signal input
flabel metal2 s 32872 200 33096 800 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 271 nsew signal input
flabel metal2 s 46984 59200 47208 59800 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 272 nsew signal input
flabel metal3 s 59200 59080 59800 59304 0 FreeSans 896 0 0 0 wbs_dat_i[18]
port 273 nsew signal input
flabel metal2 s 10696 59200 10920 59800 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 274 nsew signal input
flabel metal2 s 8680 200 8904 800 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 275 nsew signal input
flabel metal3 s 59200 32200 59800 32424 0 FreeSans 896 0 0 0 wbs_dat_i[20]
port 276 nsew signal input
flabel metal3 s 59200 57736 59800 57960 0 FreeSans 896 0 0 0 wbs_dat_i[21]
port 277 nsew signal input
flabel metal3 s 200 43624 800 43848 0 FreeSans 896 0 0 0 wbs_dat_i[22]
port 278 nsew signal input
flabel metal3 s 59200 42280 59800 42504 0 FreeSans 896 0 0 0 wbs_dat_i[23]
port 279 nsew signal input
flabel metal3 s 59200 16072 59800 16296 0 FreeSans 896 0 0 0 wbs_dat_i[24]
port 280 nsew signal input
flabel metal3 s 200 22120 800 22344 0 FreeSans 896 0 0 0 wbs_dat_i[25]
port 281 nsew signal input
flabel metal2 s 55048 59200 55272 59800 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 282 nsew signal input
flabel metal2 s 20104 59200 20328 59800 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 283 nsew signal input
flabel metal2 s 18088 200 18312 800 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 284 nsew signal input
flabel metal3 s 59200 32872 59800 33096 0 FreeSans 896 0 0 0 wbs_dat_i[29]
port 285 nsew signal input
flabel metal2 s 47656 200 47880 800 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 286 nsew signal input
flabel metal3 s 59200 14728 59800 14952 0 FreeSans 896 0 0 0 wbs_dat_i[30]
port 287 nsew signal input
flabel metal3 s 200 38248 800 38472 0 FreeSans 896 0 0 0 wbs_dat_i[31]
port 288 nsew signal input
flabel metal3 s 59200 616 59800 840 0 FreeSans 896 0 0 0 wbs_dat_i[3]
port 289 nsew signal input
flabel metal2 s 9352 200 9576 800 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 290 nsew signal input
flabel metal2 s 28840 200 29064 800 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 291 nsew signal input
flabel metal3 s 59200 23464 59800 23688 0 FreeSans 896 0 0 0 wbs_dat_i[6]
port 292 nsew signal input
flabel metal2 s 51016 59200 51240 59800 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 293 nsew signal input
flabel metal3 s 59200 50344 59800 50568 0 FreeSans 896 0 0 0 wbs_dat_i[8]
port 294 nsew signal input
flabel metal3 s 59200 1288 59800 1512 0 FreeSans 896 0 0 0 wbs_dat_i[9]
port 295 nsew signal input
flabel metal3 s 200 14728 800 14952 0 FreeSans 896 0 0 0 wbs_dat_o[0]
port 296 nsew signal tristate
flabel metal3 s 59200 31528 59800 31752 0 FreeSans 896 0 0 0 wbs_dat_o[10]
port 297 nsew signal tristate
flabel metal2 s 1288 200 1512 800 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 298 nsew signal tristate
flabel metal3 s 59200 53032 59800 53256 0 FreeSans 896 0 0 0 wbs_dat_o[12]
port 299 nsew signal tristate
flabel metal2 s 48328 59200 48552 59800 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 300 nsew signal tristate
flabel metal3 s 59200 5320 59800 5544 0 FreeSans 896 0 0 0 wbs_dat_o[14]
port 301 nsew signal tristate
flabel metal2 s 46312 59200 46536 59800 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 302 nsew signal tristate
flabel metal3 s 200 20776 800 21000 0 FreeSans 896 0 0 0 wbs_dat_o[16]
port 303 nsew signal tristate
flabel metal3 s 200 16072 800 16296 0 FreeSans 896 0 0 0 wbs_dat_o[17]
port 304 nsew signal tristate
flabel metal2 s 39592 200 39816 800 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 305 nsew signal tristate
flabel metal2 s -56 200 168 800 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 306 nsew signal tristate
flabel metal2 s 46312 200 46536 800 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 307 nsew signal tristate
flabel metal3 s 200 31528 800 31752 0 FreeSans 896 0 0 0 wbs_dat_o[20]
port 308 nsew signal tristate
flabel metal3 s 200 55048 800 55272 0 FreeSans 896 0 0 0 wbs_dat_o[21]
port 309 nsew signal tristate
flabel metal2 s 18760 59200 18984 59800 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 310 nsew signal tristate
flabel metal3 s 200 22792 800 23016 0 FreeSans 896 0 0 0 wbs_dat_o[23]
port 311 nsew signal tristate
flabel metal2 s 12040 200 12264 800 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 312 nsew signal tristate
flabel metal2 s 3976 200 4200 800 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 313 nsew signal tristate
flabel metal2 s 32872 59200 33096 59800 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 314 nsew signal tristate
flabel metal2 s 19432 59200 19656 59800 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 315 nsew signal tristate
flabel metal2 s 32200 200 32424 800 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 316 nsew signal tristate
flabel metal2 s 43624 59200 43848 59800 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 317 nsew signal tristate
flabel metal3 s 59200 15400 59800 15624 0 FreeSans 896 0 0 0 wbs_dat_o[2]
port 318 nsew signal tristate
flabel metal3 s 200 40936 800 41160 0 FreeSans 896 0 0 0 wbs_dat_o[30]
port 319 nsew signal tristate
flabel metal3 s 59200 45640 59800 45864 0 FreeSans 896 0 0 0 wbs_dat_o[31]
port 320 nsew signal tristate
flabel metal2 s 12712 200 12936 800 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 321 nsew signal tristate
flabel metal2 s 22792 200 23016 800 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 322 nsew signal tristate
flabel metal3 s 200 5992 800 6216 0 FreeSans 896 0 0 0 wbs_dat_o[5]
port 323 nsew signal tristate
flabel metal3 s 59200 44296 59800 44520 0 FreeSans 896 0 0 0 wbs_dat_o[6]
port 324 nsew signal tristate
flabel metal2 s 36232 200 36456 800 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 325 nsew signal tristate
flabel metal2 s 40264 59200 40488 59800 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 326 nsew signal tristate
flabel metal2 s 38920 59200 39144 59800 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 327 nsew signal tristate
flabel metal3 s 200 56392 800 56616 0 FreeSans 896 0 0 0 wbs_sel_i[0]
port 328 nsew signal input
flabel metal2 s 5992 59200 6216 59800 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 329 nsew signal input
flabel metal2 s 43624 200 43848 800 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 330 nsew signal input
flabel metal3 s 200 13384 800 13608 0 FreeSans 896 0 0 0 wbs_sel_i[3]
port 331 nsew signal input
flabel metal3 s 200 49672 800 49896 0 FreeSans 896 0 0 0 wbs_stb_i
port 332 nsew signal input
flabel metal3 s 59200 29512 59800 29736 0 FreeSans 896 0 0 0 wbs_we_i
port 333 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 43288 48328 43288 48328 0 _000_
rlabel metal2 44296 49000 44296 49000 0 _001_
rlabel metal2 47656 48328 47656 48328 0 _002_
rlabel metal3 45080 48888 45080 48888 0 _003_
rlabel metal2 48664 50400 48664 50400 0 _004_
rlabel metal2 46424 50288 46424 50288 0 _005_
rlabel metal3 48888 51576 48888 51576 0 _006_
rlabel metal2 46760 51744 46760 51744 0 _007_
rlabel metal2 45528 49280 45528 49280 0 _008_
rlabel metal2 44744 48552 44744 48552 0 _009_
rlabel metal3 49224 37464 49224 37464 0 _010_
rlabel metal3 45304 51352 45304 51352 0 _011_
rlabel metal2 44520 51800 44520 51800 0 _012_
rlabel metal2 44856 52584 44856 52584 0 _013_
rlabel metal2 45640 51632 45640 51632 0 _014_
rlabel metal3 45192 52920 45192 52920 0 _015_
rlabel metal3 44856 53144 44856 53144 0 _016_
rlabel metal3 45304 49784 45304 49784 0 _017_
rlabel metal2 44184 51464 44184 51464 0 _018_
rlabel metal3 48328 53704 48328 53704 0 _019_
rlabel metal2 48216 50120 48216 50120 0 _020_
rlabel metal2 54488 47936 54488 47936 0 _021_
rlabel metal2 54600 47152 54600 47152 0 _022_
rlabel metal2 52248 49784 52248 49784 0 _023_
rlabel metal3 53760 48776 53760 48776 0 _024_
rlabel metal2 53648 49224 53648 49224 0 _025_
rlabel metal2 51800 48720 51800 48720 0 _026_
rlabel metal2 51968 48216 51968 48216 0 _027_
rlabel metal3 53200 49000 53200 49000 0 _028_
rlabel metal3 52640 50008 52640 50008 0 _029_
rlabel metal2 51408 52024 51408 52024 0 _030_
rlabel metal2 50008 39984 50008 39984 0 _031_
rlabel metal2 51576 47208 51576 47208 0 _032_
rlabel metal2 51016 42168 51016 42168 0 _033_
rlabel metal2 52416 46760 52416 46760 0 _034_
rlabel metal2 52136 45752 52136 45752 0 _035_
rlabel metal3 50792 46424 50792 46424 0 _036_
rlabel metal3 51856 45864 51856 45864 0 _037_
rlabel metal2 52024 46312 52024 46312 0 _038_
rlabel metal2 52640 43848 52640 43848 0 _039_
rlabel metal2 52808 40936 52808 40936 0 _040_
rlabel metal2 49784 38976 49784 38976 0 _041_
rlabel metal3 53648 41384 53648 41384 0 _042_
rlabel metal3 54208 41720 54208 41720 0 _043_
rlabel metal3 53144 41832 53144 41832 0 _044_
rlabel metal3 52696 41944 52696 41944 0 _045_
rlabel metal2 53816 44240 53816 44240 0 _046_
rlabel metal2 52640 46648 52640 46648 0 _047_
rlabel metal2 53480 46424 53480 46424 0 _048_
rlabel metal2 53368 45808 53368 45808 0 _049_
rlabel metal2 48440 42000 48440 42000 0 _050_
rlabel metal2 49112 41720 49112 41720 0 _051_
rlabel metal3 49000 42840 49000 42840 0 _052_
rlabel metal3 49112 41832 49112 41832 0 _053_
rlabel metal3 47040 44968 47040 44968 0 _054_
rlabel metal2 47208 46032 47208 46032 0 _055_
rlabel metal2 47600 45864 47600 45864 0 _056_
rlabel metal2 48216 44800 48216 44800 0 _057_
rlabel metal2 47768 45360 47768 45360 0 _058_
rlabel metal3 47208 44856 47208 44856 0 _059_
rlabel metal3 50512 44184 50512 44184 0 _060_
rlabel metal2 55272 45920 55272 45920 0 _061_
rlabel metal2 47880 47264 47880 47264 0 _062_
rlabel metal2 47544 49504 47544 49504 0 _063_
rlabel metal3 47936 48328 47936 48328 0 _064_
rlabel metal2 48160 47432 48160 47432 0 _065_
rlabel metal2 47096 46032 47096 46032 0 _066_
rlabel metal2 53088 44296 53088 44296 0 _067_
rlabel metal2 53928 44352 53928 44352 0 _068_
rlabel metal2 45080 44520 45080 44520 0 _069_
rlabel metal3 45304 44296 45304 44296 0 _070_
rlabel via2 48104 41944 48104 41944 0 _071_
rlabel metal3 47824 41048 47824 41048 0 _072_
rlabel metal2 46760 41272 46760 41272 0 _073_
rlabel metal3 46984 41160 46984 41160 0 _074_
rlabel metal2 46032 44520 46032 44520 0 _075_
rlabel metal2 45640 44576 45640 44576 0 _076_
rlabel metal2 43736 44800 43736 44800 0 _077_
rlabel metal2 42840 45360 42840 45360 0 _078_
rlabel metal3 42448 26264 42448 26264 0 _079_
rlabel metal2 43400 45136 43400 45136 0 _080_
rlabel metal2 42392 47096 42392 47096 0 _081_
rlabel metal2 46312 45472 46312 45472 0 _082_
rlabel metal3 45360 47208 45360 47208 0 _083_
rlabel metal3 47040 41384 47040 41384 0 _084_
rlabel metal2 45864 47544 45864 47544 0 _085_
rlabel metal2 47936 49784 47936 49784 0 _086_
rlabel metal2 48104 52024 48104 52024 0 _087_
rlabel metal2 48216 51576 48216 51576 0 _088_
rlabel metal2 47656 50904 47656 50904 0 _089_
rlabel via2 46536 49000 46536 49000 0 _090_
rlabel metal3 47040 48216 47040 48216 0 _091_
rlabel metal2 44408 47488 44408 47488 0 _092_
rlabel metal2 42616 48496 42616 48496 0 _093_
rlabel metal2 41720 48384 41720 48384 0 _094_
rlabel metal3 58338 37128 58338 37128 0 io_in[0]
rlabel metal2 55384 47600 55384 47600 0 io_in[1]
rlabel metal2 5824 55384 5824 55384 0 io_in[2]
rlabel metal3 54544 55384 54544 55384 0 io_in[3]
rlabel metal2 28560 3416 28560 3416 0 io_in[4]
rlabel metal3 58338 23016 58338 23016 0 io_in[5]
rlabel metal2 45584 56280 45584 56280 0 io_in[6]
rlabel metal3 57680 55160 57680 55160 0 io_in[7]
rlabel metal2 57400 19768 57400 19768 0 io_in[8]
rlabel metal2 11592 2086 11592 2086 0 io_in[9]
rlabel metal3 1358 53256 1358 53256 0 io_out[0]
rlabel metal2 56056 40712 56056 40712 0 io_out[1]
rlabel metal3 1358 54600 1358 54600 0 io_out[2]
rlabel metal2 49224 2086 49224 2086 0 io_out[3]
rlabel metal3 57330 49672 57330 49672 0 io_out[4]
rlabel metal3 1358 25032 1358 25032 0 io_out[5]
rlabel metal2 2968 56168 2968 56168 0 io_out[6]
rlabel metal2 55384 35336 55384 35336 0 io_out[7]
rlabel metal2 57400 56280 57400 56280 0 io_out[8]
rlabel metal2 12040 57610 12040 57610 0 io_out[9]
rlabel metal2 55608 37520 55608 37520 0 net1
rlabel metal3 26880 3640 26880 3640 0 net10
rlabel metal2 29792 56280 29792 56280 0 net100
rlabel metal2 33824 56280 33824 56280 0 net101
rlabel metal2 58072 13720 58072 13720 0 net102
rlabel metal3 1302 14952 1302 14952 0 net103
rlabel metal2 46536 2030 46536 2030 0 net104
rlabel metal2 58072 15736 58072 15736 0 net105
rlabel metal2 12936 2030 12936 2030 0 net106
rlabel metal2 23016 2030 23016 2030 0 net107
rlabel metal3 1302 6216 1302 6216 0 net108
rlabel metal2 58072 44856 58072 44856 0 net109
rlabel metal2 55160 6300 55160 6300 0 net11
rlabel metal2 36456 2030 36456 2030 0 net110
rlabel metal2 41048 56504 41048 56504 0 net111
rlabel metal2 39200 56280 39200 56280 0 net112
rlabel metal3 58674 31528 58674 31528 0 net113
rlabel metal2 1512 2030 1512 2030 0 net114
rlabel metal2 58072 53368 58072 53368 0 net115
rlabel metal2 48720 56280 48720 56280 0 net116
rlabel metal2 58072 5768 58072 5768 0 net117
rlabel metal3 47264 56280 47264 56280 0 net118
rlabel metal3 1302 21000 1302 21000 0 net119
rlabel metal2 3528 52752 3528 52752 0 net12
rlabel metal3 1302 16296 1302 16296 0 net120
rlabel metal2 39816 2030 39816 2030 0 net121
rlabel metal2 168 1190 168 1190 0 net122
rlabel metal3 1302 31528 1302 31528 0 net123
rlabel metal3 1302 55272 1302 55272 0 net124
rlabel metal2 19040 56280 19040 56280 0 net125
rlabel metal3 1302 23016 1302 23016 0 net126
rlabel metal2 12264 2590 12264 2590 0 net127
rlabel metal2 4200 2030 4200 2030 0 net128
rlabel metal2 33152 56280 33152 56280 0 net129
rlabel metal2 55160 40824 55160 40824 0 net13
rlabel metal2 19712 56280 19712 56280 0 net130
rlabel metal2 32424 1246 32424 1246 0 net131
rlabel metal2 43904 56280 43904 56280 0 net132
rlabel metal3 1638 40936 1638 40936 0 net133
rlabel metal3 58674 45640 58674 45640 0 net134
rlabel metal2 3752 53592 3752 53592 0 net14
rlabel metal2 50624 4536 50624 4536 0 net15
rlabel metal3 57120 49112 57120 49112 0 net16
rlabel metal2 3080 25368 3080 25368 0 net17
rlabel metal2 4536 56056 4536 56056 0 net18
rlabel metal3 57120 35000 57120 35000 0 net19
rlabel metal3 56840 47544 56840 47544 0 net2
rlabel metal1 56392 54264 56392 54264 0 net20
rlabel metal3 28336 54376 28336 54376 0 net21
rlabel metal2 48888 54880 48888 54880 0 net22
rlabel metal2 55272 48944 55272 48944 0 net23
rlabel metal3 45752 25592 45752 25592 0 net24
rlabel metal2 58072 52808 58072 52808 0 net25
rlabel metal2 22400 56280 22400 56280 0 net26
rlabel metal3 1358 2184 1358 2184 0 net27
rlabel metal3 1302 14280 1302 14280 0 net28
rlabel metal3 1302 39816 1302 39816 0 net29
rlabel metal2 47992 53536 47992 53536 0 net3
rlabel metal2 39144 2030 39144 2030 0 net30
rlabel metal2 4872 57778 4872 57778 0 net31
rlabel metal3 36792 56280 36792 56280 0 net32
rlabel metal2 35112 2030 35112 2030 0 net33
rlabel metal3 1302 12712 1302 12712 0 net34
rlabel metal2 58128 4872 58128 4872 0 net35
rlabel metal3 1302 28392 1302 28392 0 net36
rlabel metal2 16296 2030 16296 2030 0 net37
rlabel metal3 1638 31080 1638 31080 0 net38
rlabel metal2 58072 11032 58072 11032 0 net39
rlabel metal3 56616 55944 56616 55944 0 net4
rlabel metal3 1302 39144 1302 39144 0 net40
rlabel metal2 55944 2744 55944 2744 0 net41
rlabel metal2 27104 56280 27104 56280 0 net42
rlabel metal2 11032 57792 11032 57792 0 net43
rlabel metal3 1302 52584 1302 52584 0 net44
rlabel metal2 57960 57218 57960 57218 0 net45
rlabel metal2 1848 26880 1848 26880 0 net46
rlabel metal3 1246 21672 1246 21672 0 net47
rlabel metal2 14952 2030 14952 2030 0 net48
rlabel metal2 57960 2030 57960 2030 0 net49
rlabel metal2 30744 3696 30744 3696 0 net5
rlabel metal3 1638 45640 1638 45640 0 net50
rlabel metal2 58072 3976 58072 3976 0 net51
rlabel metal3 1302 44520 1302 44520 0 net52
rlabel metal2 47208 2030 47208 2030 0 net53
rlabel metal2 22344 2030 22344 2030 0 net54
rlabel metal3 1302 35112 1302 35112 0 net55
rlabel metal2 28392 57778 28392 57778 0 net56
rlabel metal2 3584 55160 3584 55160 0 net57
rlabel metal3 58674 28392 58674 28392 0 net58
rlabel metal2 55944 1246 55944 1246 0 net59
rlabel metal2 55160 23072 55160 23072 0 net6
rlabel metal2 38528 56280 38528 56280 0 net60
rlabel metal2 48216 3304 48216 3304 0 net61
rlabel metal3 2016 54712 2016 54712 0 net62
rlabel metal2 14336 56280 14336 56280 0 net63
rlabel metal2 49560 57792 49560 57792 0 net64
rlabel metal2 16352 56280 16352 56280 0 net65
rlabel metal2 58072 30744 58072 30744 0 net66
rlabel metal2 9632 56280 9632 56280 0 net67
rlabel metal3 58674 40488 58674 40488 0 net68
rlabel metal3 1974 58408 1974 58408 0 net69
rlabel metal3 46760 55944 46760 55944 0 net7
rlabel metal3 1302 47208 1302 47208 0 net70
rlabel metal2 58072 46648 58072 46648 0 net71
rlabel metal2 58072 51352 58072 51352 0 net72
rlabel metal3 1302 19656 1302 19656 0 net73
rlabel metal2 51240 798 51240 798 0 net74
rlabel metal2 57456 55160 57456 55160 0 net75
rlabel metal3 1302 51240 1302 51240 0 net76
rlabel metal2 58072 24584 58072 24584 0 net77
rlabel metal3 1302 53928 1302 53928 0 net78
rlabel metal2 18984 2030 18984 2030 0 net79
rlabel metal2 55160 53816 55160 53816 0 net8
rlabel metal3 1302 4872 1302 4872 0 net80
rlabel metal2 58072 39256 58072 39256 0 net81
rlabel metal2 13664 56280 13664 56280 0 net82
rlabel metal3 58912 57400 58912 57400 0 net83
rlabel metal3 1302 18312 1302 18312 0 net84
rlabel metal2 31808 56280 31808 56280 0 net85
rlabel metal2 3528 2030 3528 2030 0 net86
rlabel metal2 50568 1246 50568 1246 0 net87
rlabel metal3 1246 45192 1246 45192 0 net88
rlabel metal2 4312 55300 4312 55300 0 net89
rlabel metal2 54880 20160 54880 20160 0 net9
rlabel metal2 24360 2030 24360 2030 0 net90
rlabel metal2 41720 56448 41720 56448 0 net91
rlabel metal2 58072 48104 58072 48104 0 net92
rlabel metal3 13328 55160 13328 55160 0 net93
rlabel metal2 57400 31304 57400 31304 0 net94
rlabel metal3 1302 10248 1302 10248 0 net95
rlabel metal3 1302 9576 1302 9576 0 net96
rlabel metal2 37800 56448 37800 56448 0 net97
rlabel metal2 21392 56280 21392 56280 0 net98
rlabel metal3 1246 40488 1246 40488 0 net99
rlabel metal2 57288 45920 57288 45920 0 top_wrapper.A1
rlabel metal2 51688 52416 51688 52416 0 top_wrapper.E1
rlabel metal2 48328 36904 48328 36904 0 top_wrapper.H1
rlabel metal2 55888 46872 55888 46872 0 top_wrapper.H2
rlabel metal2 42616 25984 42616 25984 0 top_wrapper.I1
rlabel metal2 41384 49672 41384 49672 0 top_wrapper.I2
rlabel metal2 54376 36568 54376 36568 0 top_wrapper.J1
rlabel metal3 52920 54600 52920 54600 0 top_wrapper.J2
rlabel metal2 44296 53760 44296 53760 0 top_wrapper.J3
rlabel metal2 41944 51856 41944 51856 0 top_wrapper.M00
rlabel metal2 49896 48720 49896 48720 0 top_wrapper.in1C\[0\]
rlabel metal3 50736 48104 50736 48104 0 top_wrapper.in1C\[1\]
rlabel metal2 50456 50456 50456 50456 0 top_wrapper.in1C\[2\]
rlabel metal2 52808 48552 52808 48552 0 top_wrapper.in1C\[3\]
rlabel metal2 49280 45640 49280 45640 0 top_wrapper.in1C\[4\]
rlabel metal2 48776 45640 48776 45640 0 top_wrapper.in2C\[0\]
rlabel metal3 49728 50344 49728 50344 0 top_wrapper.in2C\[1\]
rlabel metal2 53480 51912 53480 51912 0 top_wrapper.in2C\[2\]
rlabel metal2 48888 50008 48888 50008 0 top_wrapper.in2C\[3\]
rlabel metal3 45024 50456 45024 50456 0 top_wrapper.in2C\[4\]
rlabel metal3 58338 4200 58338 4200 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
