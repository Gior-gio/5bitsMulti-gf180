magic
tech gf180mcuC
magscale 1 5
timestamp 1670119372
<< obsm1 >>
rect 672 855 29288 28377
<< metal2 >>
rect 308 29600 420 29900
rect 644 29600 756 29900
rect 980 29600 1092 29900
rect 1316 29600 1428 29900
rect 1652 29600 1764 29900
rect 1988 29600 2100 29900
rect 2324 29600 2436 29900
rect 2660 29600 2772 29900
rect 2996 29600 3108 29900
rect 3332 29600 3444 29900
rect 3668 29600 3780 29900
rect 4340 29600 4452 29900
rect 4676 29600 4788 29900
rect 5012 29600 5124 29900
rect 5348 29600 5460 29900
rect 5684 29600 5796 29900
rect 6020 29600 6132 29900
rect 6356 29600 6468 29900
rect 6692 29600 6804 29900
rect 7028 29600 7140 29900
rect 7364 29600 7476 29900
rect 7700 29600 7812 29900
rect 8036 29600 8148 29900
rect 8708 29600 8820 29900
rect 9044 29600 9156 29900
rect 9380 29600 9492 29900
rect 9716 29600 9828 29900
rect 10052 29600 10164 29900
rect 10388 29600 10500 29900
rect 10724 29600 10836 29900
rect 11060 29600 11172 29900
rect 11396 29600 11508 29900
rect 11732 29600 11844 29900
rect 12068 29600 12180 29900
rect 12404 29600 12516 29900
rect 13076 29600 13188 29900
rect 13412 29600 13524 29900
rect 13748 29600 13860 29900
rect 14084 29600 14196 29900
rect 14420 29600 14532 29900
rect 14756 29600 14868 29900
rect 15092 29600 15204 29900
rect 15428 29600 15540 29900
rect 15764 29600 15876 29900
rect 16100 29600 16212 29900
rect 16436 29600 16548 29900
rect 16772 29600 16884 29900
rect 17444 29600 17556 29900
rect 17780 29600 17892 29900
rect 18116 29600 18228 29900
rect 18452 29600 18564 29900
rect 18788 29600 18900 29900
rect 19124 29600 19236 29900
rect 19460 29600 19572 29900
rect 19796 29600 19908 29900
rect 20132 29600 20244 29900
rect 20468 29600 20580 29900
rect 20804 29600 20916 29900
rect 21140 29600 21252 29900
rect 21812 29600 21924 29900
rect 22148 29600 22260 29900
rect 22484 29600 22596 29900
rect 22820 29600 22932 29900
rect 23156 29600 23268 29900
rect 23492 29600 23604 29900
rect 23828 29600 23940 29900
rect 24164 29600 24276 29900
rect 24500 29600 24612 29900
rect 24836 29600 24948 29900
rect 25172 29600 25284 29900
rect 25508 29600 25620 29900
rect 26180 29600 26292 29900
rect 26516 29600 26628 29900
rect 26852 29600 26964 29900
rect 27188 29600 27300 29900
rect 27524 29600 27636 29900
rect 27860 29600 27972 29900
rect 28196 29600 28308 29900
rect 28532 29600 28644 29900
rect 28868 29600 28980 29900
rect 29204 29600 29316 29900
rect 29540 29600 29652 29900
rect 29876 29600 29988 29900
rect -28 100 84 400
rect 308 100 420 400
rect 644 100 756 400
rect 980 100 1092 400
rect 1316 100 1428 400
rect 1652 100 1764 400
rect 1988 100 2100 400
rect 2324 100 2436 400
rect 2660 100 2772 400
rect 2996 100 3108 400
rect 3332 100 3444 400
rect 3668 100 3780 400
rect 4340 100 4452 400
rect 4676 100 4788 400
rect 5012 100 5124 400
rect 5348 100 5460 400
rect 5684 100 5796 400
rect 6020 100 6132 400
rect 6356 100 6468 400
rect 6692 100 6804 400
rect 7028 100 7140 400
rect 7364 100 7476 400
rect 7700 100 7812 400
rect 8036 100 8148 400
rect 8708 100 8820 400
rect 9044 100 9156 400
rect 9380 100 9492 400
rect 9716 100 9828 400
rect 10052 100 10164 400
rect 10388 100 10500 400
rect 10724 100 10836 400
rect 11060 100 11172 400
rect 11396 100 11508 400
rect 11732 100 11844 400
rect 12068 100 12180 400
rect 12404 100 12516 400
rect 13076 100 13188 400
rect 13412 100 13524 400
rect 13748 100 13860 400
rect 14084 100 14196 400
rect 14420 100 14532 400
rect 14756 100 14868 400
rect 15092 100 15204 400
rect 15428 100 15540 400
rect 15764 100 15876 400
rect 16100 100 16212 400
rect 16436 100 16548 400
rect 16772 100 16884 400
rect 17444 100 17556 400
rect 17780 100 17892 400
rect 18116 100 18228 400
rect 18452 100 18564 400
rect 18788 100 18900 400
rect 19124 100 19236 400
rect 19460 100 19572 400
rect 19796 100 19908 400
rect 20132 100 20244 400
rect 20468 100 20580 400
rect 20804 100 20916 400
rect 21140 100 21252 400
rect 21812 100 21924 400
rect 22148 100 22260 400
rect 22484 100 22596 400
rect 22820 100 22932 400
rect 23156 100 23268 400
rect 23492 100 23604 400
rect 23828 100 23940 400
rect 24164 100 24276 400
rect 24500 100 24612 400
rect 24836 100 24948 400
rect 25172 100 25284 400
rect 25508 100 25620 400
rect 26180 100 26292 400
rect 26516 100 26628 400
rect 26852 100 26964 400
rect 27188 100 27300 400
rect 27524 100 27636 400
rect 27860 100 27972 400
rect 28196 100 28308 400
rect 28532 100 28644 400
rect 28868 100 28980 400
rect 29204 100 29316 400
rect 29540 100 29652 400
<< obsm2 >>
rect 70 29570 278 29666
rect 450 29570 614 29666
rect 786 29570 950 29666
rect 1122 29570 1286 29666
rect 1458 29570 1622 29666
rect 1794 29570 1958 29666
rect 2130 29570 2294 29666
rect 2466 29570 2630 29666
rect 2802 29570 2966 29666
rect 3138 29570 3302 29666
rect 3474 29570 3638 29666
rect 3810 29570 4310 29666
rect 4482 29570 4646 29666
rect 4818 29570 4982 29666
rect 5154 29570 5318 29666
rect 5490 29570 5654 29666
rect 5826 29570 5990 29666
rect 6162 29570 6326 29666
rect 6498 29570 6662 29666
rect 6834 29570 6998 29666
rect 7170 29570 7334 29666
rect 7506 29570 7670 29666
rect 7842 29570 8006 29666
rect 8178 29570 8678 29666
rect 8850 29570 9014 29666
rect 9186 29570 9350 29666
rect 9522 29570 9686 29666
rect 9858 29570 10022 29666
rect 10194 29570 10358 29666
rect 10530 29570 10694 29666
rect 10866 29570 11030 29666
rect 11202 29570 11366 29666
rect 11538 29570 11702 29666
rect 11874 29570 12038 29666
rect 12210 29570 12374 29666
rect 12546 29570 13046 29666
rect 13218 29570 13382 29666
rect 13554 29570 13718 29666
rect 13890 29570 14054 29666
rect 14226 29570 14390 29666
rect 14562 29570 14726 29666
rect 14898 29570 15062 29666
rect 15234 29570 15398 29666
rect 15570 29570 15734 29666
rect 15906 29570 16070 29666
rect 16242 29570 16406 29666
rect 16578 29570 16742 29666
rect 16914 29570 17414 29666
rect 17586 29570 17750 29666
rect 17922 29570 18086 29666
rect 18258 29570 18422 29666
rect 18594 29570 18758 29666
rect 18930 29570 19094 29666
rect 19266 29570 19430 29666
rect 19602 29570 19766 29666
rect 19938 29570 20102 29666
rect 20274 29570 20438 29666
rect 20610 29570 20774 29666
rect 20946 29570 21110 29666
rect 21282 29570 21782 29666
rect 21954 29570 22118 29666
rect 22290 29570 22454 29666
rect 22626 29570 22790 29666
rect 22962 29570 23126 29666
rect 23298 29570 23462 29666
rect 23634 29570 23798 29666
rect 23970 29570 24134 29666
rect 24306 29570 24470 29666
rect 24642 29570 24806 29666
rect 24978 29570 25142 29666
rect 25314 29570 25478 29666
rect 25650 29570 26150 29666
rect 26322 29570 26486 29666
rect 26658 29570 26822 29666
rect 26994 29570 27158 29666
rect 27330 29570 27494 29666
rect 27666 29570 27830 29666
rect 28002 29570 28166 29666
rect 28338 29570 28502 29666
rect 28674 29570 28838 29666
rect 29010 29570 29174 29666
rect 29346 29570 29510 29666
rect 29682 29570 29846 29666
rect 70 430 29890 29570
rect 114 70 278 430
rect 450 70 614 430
rect 786 70 950 430
rect 1122 70 1286 430
rect 1458 70 1622 430
rect 1794 70 1958 430
rect 2130 70 2294 430
rect 2466 70 2630 430
rect 2802 70 2966 430
rect 3138 70 3302 430
rect 3474 70 3638 430
rect 3810 70 4310 430
rect 4482 70 4646 430
rect 4818 70 4982 430
rect 5154 70 5318 430
rect 5490 70 5654 430
rect 5826 70 5990 430
rect 6162 70 6326 430
rect 6498 70 6662 430
rect 6834 70 6998 430
rect 7170 70 7334 430
rect 7506 70 7670 430
rect 7842 70 8006 430
rect 8178 70 8678 430
rect 8850 70 9014 430
rect 9186 70 9350 430
rect 9522 70 9686 430
rect 9858 70 10022 430
rect 10194 70 10358 430
rect 10530 70 10694 430
rect 10866 70 11030 430
rect 11202 70 11366 430
rect 11538 70 11702 430
rect 11874 70 12038 430
rect 12210 70 12374 430
rect 12546 70 13046 430
rect 13218 70 13382 430
rect 13554 70 13718 430
rect 13890 70 14054 430
rect 14226 70 14390 430
rect 14562 70 14726 430
rect 14898 70 15062 430
rect 15234 70 15398 430
rect 15570 70 15734 430
rect 15906 70 16070 430
rect 16242 70 16406 430
rect 16578 70 16742 430
rect 16914 70 17414 430
rect 17586 70 17750 430
rect 17922 70 18086 430
rect 18258 70 18422 430
rect 18594 70 18758 430
rect 18930 70 19094 430
rect 19266 70 19430 430
rect 19602 70 19766 430
rect 19938 70 20102 430
rect 20274 70 20438 430
rect 20610 70 20774 430
rect 20946 70 21110 430
rect 21282 70 21782 430
rect 21954 70 22118 430
rect 22290 70 22454 430
rect 22626 70 22790 430
rect 22962 70 23126 430
rect 23298 70 23462 430
rect 23634 70 23798 430
rect 23970 70 24134 430
rect 24306 70 24470 430
rect 24642 70 24806 430
rect 24978 70 25142 430
rect 25314 70 25478 430
rect 25650 70 26150 430
rect 26322 70 26486 430
rect 26658 70 26822 430
rect 26994 70 27158 430
rect 27330 70 27494 430
rect 27666 70 27830 430
rect 28002 70 28166 430
rect 28338 70 28502 430
rect 28674 70 28838 430
rect 29010 70 29174 430
rect 29346 70 29510 430
rect 29682 70 29890 430
rect 70 65 29890 70
<< metal3 >>
rect 100 29876 400 29988
rect 100 29540 400 29652
rect 29600 29540 29900 29652
rect 100 29204 400 29316
rect 29600 29204 29900 29316
rect 100 28868 400 28980
rect 29600 28868 29900 28980
rect 100 28532 400 28644
rect 29600 28532 29900 28644
rect 100 28196 400 28308
rect 29600 28196 29900 28308
rect 100 27860 400 27972
rect 29600 27860 29900 27972
rect 100 27524 400 27636
rect 29600 27524 29900 27636
rect 100 27188 400 27300
rect 29600 27188 29900 27300
rect 100 26852 400 26964
rect 29600 26852 29900 26964
rect 100 26516 400 26628
rect 29600 26516 29900 26628
rect 100 26180 400 26292
rect 29600 26180 29900 26292
rect 100 25508 400 25620
rect 29600 25508 29900 25620
rect 100 25172 400 25284
rect 29600 25172 29900 25284
rect 100 24836 400 24948
rect 29600 24836 29900 24948
rect 100 24500 400 24612
rect 29600 24500 29900 24612
rect 100 24164 400 24276
rect 29600 24164 29900 24276
rect 100 23828 400 23940
rect 29600 23828 29900 23940
rect 100 23492 400 23604
rect 29600 23492 29900 23604
rect 100 23156 400 23268
rect 29600 23156 29900 23268
rect 100 22820 400 22932
rect 29600 22820 29900 22932
rect 100 22484 400 22596
rect 29600 22484 29900 22596
rect 100 22148 400 22260
rect 29600 22148 29900 22260
rect 100 21812 400 21924
rect 29600 21812 29900 21924
rect 100 21140 400 21252
rect 29600 21140 29900 21252
rect 100 20804 400 20916
rect 29600 20804 29900 20916
rect 100 20468 400 20580
rect 29600 20468 29900 20580
rect 100 20132 400 20244
rect 29600 20132 29900 20244
rect 100 19796 400 19908
rect 29600 19796 29900 19908
rect 100 19460 400 19572
rect 29600 19460 29900 19572
rect 100 19124 400 19236
rect 29600 19124 29900 19236
rect 100 18788 400 18900
rect 29600 18788 29900 18900
rect 100 18452 400 18564
rect 29600 18452 29900 18564
rect 100 18116 400 18228
rect 29600 18116 29900 18228
rect 100 17780 400 17892
rect 29600 17780 29900 17892
rect 100 17444 400 17556
rect 29600 17444 29900 17556
rect 100 16772 400 16884
rect 29600 16772 29900 16884
rect 100 16436 400 16548
rect 29600 16436 29900 16548
rect 100 16100 400 16212
rect 29600 16100 29900 16212
rect 100 15764 400 15876
rect 29600 15764 29900 15876
rect 100 15428 400 15540
rect 29600 15428 29900 15540
rect 100 15092 400 15204
rect 29600 15092 29900 15204
rect 100 14756 400 14868
rect 29600 14756 29900 14868
rect 100 14420 400 14532
rect 29600 14420 29900 14532
rect 100 14084 400 14196
rect 29600 14084 29900 14196
rect 100 13748 400 13860
rect 29600 13748 29900 13860
rect 100 13412 400 13524
rect 29600 13412 29900 13524
rect 100 13076 400 13188
rect 29600 13076 29900 13188
rect 100 12404 400 12516
rect 29600 12404 29900 12516
rect 100 12068 400 12180
rect 29600 12068 29900 12180
rect 100 11732 400 11844
rect 29600 11732 29900 11844
rect 100 11396 400 11508
rect 29600 11396 29900 11508
rect 100 11060 400 11172
rect 29600 11060 29900 11172
rect 100 10724 400 10836
rect 29600 10724 29900 10836
rect 100 10388 400 10500
rect 29600 10388 29900 10500
rect 100 10052 400 10164
rect 29600 10052 29900 10164
rect 100 9716 400 9828
rect 29600 9716 29900 9828
rect 100 9380 400 9492
rect 29600 9380 29900 9492
rect 100 9044 400 9156
rect 29600 9044 29900 9156
rect 100 8708 400 8820
rect 29600 8708 29900 8820
rect 100 8036 400 8148
rect 29600 8036 29900 8148
rect 100 7700 400 7812
rect 29600 7700 29900 7812
rect 100 7364 400 7476
rect 29600 7364 29900 7476
rect 100 7028 400 7140
rect 29600 7028 29900 7140
rect 100 6692 400 6804
rect 29600 6692 29900 6804
rect 100 6356 400 6468
rect 29600 6356 29900 6468
rect 100 6020 400 6132
rect 29600 6020 29900 6132
rect 100 5684 400 5796
rect 29600 5684 29900 5796
rect 100 5348 400 5460
rect 29600 5348 29900 5460
rect 100 5012 400 5124
rect 29600 5012 29900 5124
rect 100 4676 400 4788
rect 29600 4676 29900 4788
rect 100 4340 400 4452
rect 29600 4340 29900 4452
rect 100 3668 400 3780
rect 29600 3668 29900 3780
rect 100 3332 400 3444
rect 29600 3332 29900 3444
rect 100 2996 400 3108
rect 29600 2996 29900 3108
rect 100 2660 400 2772
rect 29600 2660 29900 2772
rect 100 2324 400 2436
rect 29600 2324 29900 2436
rect 100 1988 400 2100
rect 29600 1988 29900 2100
rect 100 1652 400 1764
rect 29600 1652 29900 1764
rect 100 1316 400 1428
rect 29600 1316 29900 1428
rect 100 980 400 1092
rect 29600 980 29900 1092
rect 100 644 400 756
rect 29600 644 29900 756
rect 100 308 400 420
rect 29600 308 29900 420
rect 29600 -28 29900 84
<< obsm3 >>
rect 65 29174 70 29218
rect 430 29174 29570 29218
rect 65 29010 29895 29174
rect 65 28838 70 29010
rect 430 28838 29570 29010
rect 65 28674 29895 28838
rect 65 28502 70 28674
rect 430 28502 29570 28674
rect 65 28338 29895 28502
rect 65 28166 70 28338
rect 430 28166 29570 28338
rect 65 28002 29895 28166
rect 65 27830 70 28002
rect 430 27830 29570 28002
rect 65 27666 29895 27830
rect 65 27494 70 27666
rect 430 27494 29570 27666
rect 65 27330 29895 27494
rect 65 27158 70 27330
rect 430 27158 29570 27330
rect 65 26994 29895 27158
rect 65 26822 70 26994
rect 430 26822 29570 26994
rect 65 26658 29895 26822
rect 65 26486 70 26658
rect 430 26486 29570 26658
rect 65 26322 29895 26486
rect 65 26150 70 26322
rect 430 26150 29570 26322
rect 65 25650 29895 26150
rect 65 25478 70 25650
rect 430 25478 29570 25650
rect 65 25314 29895 25478
rect 65 25142 70 25314
rect 430 25142 29570 25314
rect 65 24978 29895 25142
rect 65 24806 70 24978
rect 430 24806 29570 24978
rect 65 24642 29895 24806
rect 65 24470 70 24642
rect 430 24470 29570 24642
rect 65 24306 29895 24470
rect 65 24134 70 24306
rect 430 24134 29570 24306
rect 65 23970 29895 24134
rect 65 23798 70 23970
rect 430 23798 29570 23970
rect 65 23634 29895 23798
rect 65 23462 70 23634
rect 430 23462 29570 23634
rect 65 23298 29895 23462
rect 65 23126 70 23298
rect 430 23126 29570 23298
rect 65 22962 29895 23126
rect 65 22790 70 22962
rect 430 22790 29570 22962
rect 65 22626 29895 22790
rect 65 22454 70 22626
rect 430 22454 29570 22626
rect 65 22290 29895 22454
rect 65 22118 70 22290
rect 430 22118 29570 22290
rect 65 21954 29895 22118
rect 65 21782 70 21954
rect 430 21782 29570 21954
rect 65 21282 29895 21782
rect 65 21110 70 21282
rect 430 21110 29570 21282
rect 65 20946 29895 21110
rect 65 20774 70 20946
rect 430 20774 29570 20946
rect 65 20610 29895 20774
rect 65 20438 70 20610
rect 430 20438 29570 20610
rect 65 20274 29895 20438
rect 65 20102 70 20274
rect 430 20102 29570 20274
rect 65 19938 29895 20102
rect 65 19766 70 19938
rect 430 19766 29570 19938
rect 65 19602 29895 19766
rect 65 19430 70 19602
rect 430 19430 29570 19602
rect 65 19266 29895 19430
rect 65 19094 70 19266
rect 430 19094 29570 19266
rect 65 18930 29895 19094
rect 65 18758 70 18930
rect 430 18758 29570 18930
rect 65 18594 29895 18758
rect 65 18422 70 18594
rect 430 18422 29570 18594
rect 65 18258 29895 18422
rect 65 18086 70 18258
rect 430 18086 29570 18258
rect 65 17922 29895 18086
rect 65 17750 70 17922
rect 430 17750 29570 17922
rect 65 17586 29895 17750
rect 65 17414 70 17586
rect 430 17414 29570 17586
rect 65 16914 29895 17414
rect 65 16742 70 16914
rect 430 16742 29570 16914
rect 65 16578 29895 16742
rect 65 16406 70 16578
rect 430 16406 29570 16578
rect 65 16242 29895 16406
rect 65 16070 70 16242
rect 430 16070 29570 16242
rect 65 15906 29895 16070
rect 65 15734 70 15906
rect 430 15734 29570 15906
rect 65 15570 29895 15734
rect 65 15398 70 15570
rect 430 15398 29570 15570
rect 65 15234 29895 15398
rect 65 15062 70 15234
rect 430 15062 29570 15234
rect 65 14898 29895 15062
rect 65 14726 70 14898
rect 430 14726 29570 14898
rect 65 14562 29895 14726
rect 65 14390 70 14562
rect 430 14390 29570 14562
rect 65 14226 29895 14390
rect 65 14054 70 14226
rect 430 14054 29570 14226
rect 65 13890 29895 14054
rect 65 13718 70 13890
rect 430 13718 29570 13890
rect 65 13554 29895 13718
rect 65 13382 70 13554
rect 430 13382 29570 13554
rect 65 13218 29895 13382
rect 65 13046 70 13218
rect 430 13046 29570 13218
rect 65 12546 29895 13046
rect 65 12374 70 12546
rect 430 12374 29570 12546
rect 65 12210 29895 12374
rect 65 12038 70 12210
rect 430 12038 29570 12210
rect 65 11874 29895 12038
rect 65 11702 70 11874
rect 430 11702 29570 11874
rect 65 11538 29895 11702
rect 65 11366 70 11538
rect 430 11366 29570 11538
rect 65 11202 29895 11366
rect 65 11030 70 11202
rect 430 11030 29570 11202
rect 65 10866 29895 11030
rect 65 10694 70 10866
rect 430 10694 29570 10866
rect 65 10530 29895 10694
rect 65 10358 70 10530
rect 430 10358 29570 10530
rect 65 10194 29895 10358
rect 65 10022 70 10194
rect 430 10022 29570 10194
rect 65 9858 29895 10022
rect 65 9686 70 9858
rect 430 9686 29570 9858
rect 65 9522 29895 9686
rect 65 9350 70 9522
rect 430 9350 29570 9522
rect 65 9186 29895 9350
rect 65 9014 70 9186
rect 430 9014 29570 9186
rect 65 8850 29895 9014
rect 65 8678 70 8850
rect 430 8678 29570 8850
rect 65 8178 29895 8678
rect 65 8006 70 8178
rect 430 8006 29570 8178
rect 65 7842 29895 8006
rect 65 7670 70 7842
rect 430 7670 29570 7842
rect 65 7506 29895 7670
rect 65 7334 70 7506
rect 430 7334 29570 7506
rect 65 7170 29895 7334
rect 65 6998 70 7170
rect 430 6998 29570 7170
rect 65 6834 29895 6998
rect 65 6662 70 6834
rect 430 6662 29570 6834
rect 65 6498 29895 6662
rect 65 6326 70 6498
rect 430 6326 29570 6498
rect 65 6162 29895 6326
rect 65 5990 70 6162
rect 430 5990 29570 6162
rect 65 5826 29895 5990
rect 65 5654 70 5826
rect 430 5654 29570 5826
rect 65 5490 29895 5654
rect 65 5318 70 5490
rect 430 5318 29570 5490
rect 65 5154 29895 5318
rect 65 4982 70 5154
rect 430 4982 29570 5154
rect 65 4818 29895 4982
rect 65 4646 70 4818
rect 430 4646 29570 4818
rect 65 4482 29895 4646
rect 65 4310 70 4482
rect 430 4310 29570 4482
rect 65 3810 29895 4310
rect 65 3638 70 3810
rect 430 3638 29570 3810
rect 65 3474 29895 3638
rect 65 3302 70 3474
rect 430 3302 29570 3474
rect 65 3138 29895 3302
rect 65 2966 70 3138
rect 430 2966 29570 3138
rect 65 2802 29895 2966
rect 65 2630 70 2802
rect 430 2630 29570 2802
rect 65 2466 29895 2630
rect 65 2294 70 2466
rect 430 2294 29570 2466
rect 65 2130 29895 2294
rect 65 1958 70 2130
rect 430 1958 29570 2130
rect 65 1794 29895 1958
rect 65 1622 70 1794
rect 430 1622 29570 1794
rect 65 1458 29895 1622
rect 65 1286 70 1458
rect 430 1286 29570 1458
rect 65 1122 29895 1286
rect 65 950 70 1122
rect 430 950 29570 1122
rect 65 786 29895 950
rect 65 614 70 786
rect 430 614 29570 786
rect 65 450 29895 614
rect 65 278 70 450
rect 430 278 29570 450
rect 65 114 29895 278
rect 65 70 29570 114
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< obsm4 >>
rect 26390 24313 26418 25247
<< labels >>
rlabel metal3 s 29600 18452 29900 18564 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 29600 24164 29900 24276 6 io_in[1]
port 2 nsew signal input
rlabel metal2 s 2660 29600 2772 29900 6 io_in[2]
port 3 nsew signal input
rlabel metal2 s 29204 29600 29316 29900 6 io_in[3]
port 4 nsew signal input
rlabel metal2 s 14084 100 14196 400 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 29600 11396 29900 11508 6 io_in[5]
port 6 nsew signal input
rlabel metal2 s 22820 29600 22932 29900 6 io_in[6]
port 7 nsew signal input
rlabel metal2 s 29540 29600 29652 29900 6 io_in[7]
port 8 nsew signal input
rlabel metal3 s 29600 9716 29900 9828 6 io_in[8]
port 9 nsew signal input
rlabel metal2 s 5684 100 5796 400 6 io_in[9]
port 10 nsew signal input
rlabel metal3 s 29600 26180 29900 26292 6 io_oeb[0]
port 11 nsew signal output
rlabel metal2 s 11060 29600 11172 29900 6 io_oeb[1]
port 12 nsew signal output
rlabel metal3 s 100 980 400 1092 6 io_oeb[2]
port 13 nsew signal output
rlabel metal3 s 100 7028 400 7140 6 io_oeb[3]
port 14 nsew signal output
rlabel metal3 s 100 19796 400 19908 6 io_oeb[4]
port 15 nsew signal output
rlabel metal2 s 19460 100 19572 400 6 io_oeb[5]
port 16 nsew signal output
rlabel metal2 s 2324 29600 2436 29900 6 io_oeb[6]
port 17 nsew signal output
rlabel metal2 s 18116 29600 18228 29900 6 io_oeb[7]
port 18 nsew signal output
rlabel metal2 s 17444 100 17556 400 6 io_oeb[8]
port 19 nsew signal output
rlabel metal3 s 100 6356 400 6468 6 io_oeb[9]
port 20 nsew signal output
rlabel metal3 s 100 26516 400 26628 6 io_out[0]
port 21 nsew signal output
rlabel metal3 s 29600 20468 29900 20580 6 io_out[1]
port 22 nsew signal output
rlabel metal3 s 100 27188 400 27300 6 io_out[2]
port 23 nsew signal output
rlabel metal2 s 24500 100 24612 400 6 io_out[3]
port 24 nsew signal output
rlabel metal3 s 29600 24836 29900 24948 6 io_out[4]
port 25 nsew signal output
rlabel metal3 s 100 12404 400 12516 6 io_out[5]
port 26 nsew signal output
rlabel metal2 s 1316 29600 1428 29900 6 io_out[6]
port 27 nsew signal output
rlabel metal3 s 29600 17444 29900 17556 6 io_out[7]
port 28 nsew signal output
rlabel metal2 s 28196 29600 28308 29900 6 io_out[8]
port 29 nsew signal output
rlabel metal2 s 6020 29600 6132 29900 6 io_out[9]
port 30 nsew signal output
rlabel metal3 s 29600 13412 29900 13524 6 la_data_in[0]
port 31 nsew signal input
rlabel metal2 s 10388 100 10500 400 6 la_data_in[10]
port 32 nsew signal input
rlabel metal3 s 29600 2324 29900 2436 6 la_data_in[11]
port 33 nsew signal input
rlabel metal3 s 29600 11060 29900 11172 6 la_data_in[12]
port 34 nsew signal input
rlabel metal2 s 28532 29600 28644 29900 6 la_data_in[13]
port 35 nsew signal input
rlabel metal2 s 14756 100 14868 400 6 la_data_in[14]
port 36 nsew signal input
rlabel metal3 s 29600 12404 29900 12516 6 la_data_in[15]
port 37 nsew signal input
rlabel metal2 s 308 29600 420 29900 6 la_data_in[16]
port 38 nsew signal input
rlabel metal3 s 100 29540 400 29652 6 la_data_in[17]
port 39 nsew signal input
rlabel metal2 s 8708 100 8820 400 6 la_data_in[18]
port 40 nsew signal input
rlabel metal2 s 22484 100 22596 400 6 la_data_in[19]
port 41 nsew signal input
rlabel metal2 s 22484 29600 22596 29900 6 la_data_in[1]
port 42 nsew signal input
rlabel metal2 s 11396 29600 11508 29900 6 la_data_in[20]
port 43 nsew signal input
rlabel metal3 s 29600 13076 29900 13188 6 la_data_in[21]
port 44 nsew signal input
rlabel metal3 s 100 13748 400 13860 6 la_data_in[22]
port 45 nsew signal input
rlabel metal2 s 5012 29600 5124 29900 6 la_data_in[23]
port 46 nsew signal input
rlabel metal2 s 11732 100 11844 400 6 la_data_in[24]
port 47 nsew signal input
rlabel metal2 s 14420 29600 14532 29900 6 la_data_in[25]
port 48 nsew signal input
rlabel metal3 s 29600 20804 29900 20916 6 la_data_in[26]
port 49 nsew signal input
rlabel metal2 s 26516 29600 26628 29900 6 la_data_in[27]
port 50 nsew signal input
rlabel metal3 s 100 11732 400 11844 6 la_data_in[28]
port 51 nsew signal input
rlabel metal3 s 29600 3332 29900 3444 6 la_data_in[29]
port 52 nsew signal input
rlabel metal3 s 100 27860 400 27972 6 la_data_in[2]
port 53 nsew signal input
rlabel metal3 s 29600 28196 29900 28308 6 la_data_in[30]
port 54 nsew signal input
rlabel metal3 s 29600 18788 29900 18900 6 la_data_in[31]
port 55 nsew signal input
rlabel metal3 s 100 20804 400 20916 6 la_data_in[32]
port 56 nsew signal input
rlabel metal2 s 27524 100 27636 400 6 la_data_in[33]
port 57 nsew signal input
rlabel metal3 s 29600 4676 29900 4788 6 la_data_in[34]
port 58 nsew signal input
rlabel metal2 s 24836 29600 24948 29900 6 la_data_in[35]
port 59 nsew signal input
rlabel metal2 s 3668 29600 3780 29900 6 la_data_in[36]
port 60 nsew signal input
rlabel metal2 s 26180 29600 26292 29900 6 la_data_in[37]
port 61 nsew signal input
rlabel metal3 s 100 18788 400 18900 6 la_data_in[38]
port 62 nsew signal input
rlabel metal2 s 7364 29600 7476 29900 6 la_data_in[39]
port 63 nsew signal input
rlabel metal3 s 100 1316 400 1428 6 la_data_in[3]
port 64 nsew signal input
rlabel metal2 s 13076 29600 13188 29900 6 la_data_in[40]
port 65 nsew signal input
rlabel metal2 s 7700 100 7812 400 6 la_data_in[41]
port 66 nsew signal input
rlabel metal3 s 29600 5012 29900 5124 6 la_data_in[42]
port 67 nsew signal input
rlabel metal2 s 27188 29600 27300 29900 6 la_data_in[43]
port 68 nsew signal input
rlabel metal2 s 16772 100 16884 400 6 la_data_in[44]
port 69 nsew signal input
rlabel metal3 s 29600 19124 29900 19236 6 la_data_in[45]
port 70 nsew signal input
rlabel metal3 s 100 3332 400 3444 6 la_data_in[46]
port 71 nsew signal input
rlabel metal3 s 29600 2996 29900 3108 6 la_data_in[47]
port 72 nsew signal input
rlabel metal2 s 13748 100 13860 400 6 la_data_in[48]
port 73 nsew signal input
rlabel metal3 s 100 6020 400 6132 6 la_data_in[49]
port 74 nsew signal input
rlabel metal3 s 100 21140 400 21252 6 la_data_in[4]
port 75 nsew signal input
rlabel metal3 s 100 1652 400 1764 6 la_data_in[50]
port 76 nsew signal input
rlabel metal3 s 100 16100 400 16212 6 la_data_in[51]
port 77 nsew signal input
rlabel metal2 s 8708 29600 8820 29900 6 la_data_in[52]
port 78 nsew signal input
rlabel metal3 s 29600 1316 29900 1428 6 la_data_in[53]
port 79 nsew signal input
rlabel metal3 s 29600 7028 29900 7140 6 la_data_in[54]
port 80 nsew signal input
rlabel metal3 s 100 10052 400 10164 6 la_data_in[55]
port 81 nsew signal input
rlabel metal2 s 12404 100 12516 400 6 la_data_in[56]
port 82 nsew signal input
rlabel metal2 s 19124 100 19236 400 6 la_data_in[57]
port 83 nsew signal input
rlabel metal2 s 10724 29600 10836 29900 6 la_data_in[58]
port 84 nsew signal input
rlabel metal3 s 29600 27524 29900 27636 6 la_data_in[59]
port 85 nsew signal input
rlabel metal2 s 12068 29600 12180 29900 6 la_data_in[5]
port 86 nsew signal input
rlabel metal2 s 28196 100 28308 400 6 la_data_in[60]
port 87 nsew signal input
rlabel metal2 s 9716 100 9828 400 6 la_data_in[61]
port 88 nsew signal input
rlabel metal3 s 100 16772 400 16884 6 la_data_in[62]
port 89 nsew signal input
rlabel metal3 s 29600 5684 29900 5796 6 la_data_in[63]
port 90 nsew signal input
rlabel metal2 s 3668 100 3780 400 6 la_data_in[6]
port 91 nsew signal input
rlabel metal2 s 3332 29600 3444 29900 6 la_data_in[7]
port 92 nsew signal input
rlabel metal2 s 7700 29600 7812 29900 6 la_data_in[8]
port 93 nsew signal input
rlabel metal3 s 100 3668 400 3780 6 la_data_in[9]
port 94 nsew signal input
rlabel metal3 s 29600 -28 29900 84 6 la_data_out[0]
port 95 nsew signal output
rlabel metal2 s 28868 29600 28980 29900 6 la_data_out[10]
port 96 nsew signal output
rlabel metal3 s 100 13412 400 13524 6 la_data_out[11]
port 97 nsew signal output
rlabel metal3 s 100 10724 400 10836 6 la_data_out[12]
port 98 nsew signal output
rlabel metal2 s 7364 100 7476 400 6 la_data_out[13]
port 99 nsew signal output
rlabel metal2 s 28868 100 28980 400 6 la_data_out[14]
port 100 nsew signal output
rlabel metal3 s 100 22820 400 22932 6 la_data_out[15]
port 101 nsew signal output
rlabel metal3 s 29600 1652 29900 1764 6 la_data_out[16]
port 102 nsew signal output
rlabel metal3 s 100 22148 400 22260 6 la_data_out[17]
port 103 nsew signal output
rlabel metal2 s 23492 100 23604 400 6 la_data_out[18]
port 104 nsew signal output
rlabel metal2 s 11060 100 11172 400 6 la_data_out[19]
port 105 nsew signal output
rlabel metal3 s 100 14084 400 14196 6 la_data_out[1]
port 106 nsew signal output
rlabel metal3 s 100 17444 400 17556 6 la_data_out[20]
port 107 nsew signal output
rlabel metal2 s 14084 29600 14196 29900 6 la_data_out[21]
port 108 nsew signal output
rlabel metal2 s 1652 29600 1764 29900 6 la_data_out[22]
port 109 nsew signal output
rlabel metal3 s 29600 14084 29900 14196 6 la_data_out[23]
port 110 nsew signal output
rlabel metal2 s 27860 100 27972 400 6 la_data_out[24]
port 111 nsew signal output
rlabel metal2 s 19124 29600 19236 29900 6 la_data_out[25]
port 112 nsew signal output
rlabel metal2 s 24164 100 24276 400 6 la_data_out[26]
port 113 nsew signal output
rlabel metal2 s 644 29600 756 29900 6 la_data_out[27]
port 114 nsew signal output
rlabel metal2 s 7028 29600 7140 29900 6 la_data_out[28]
port 115 nsew signal output
rlabel metal2 s 24500 29600 24612 29900 6 la_data_out[29]
port 116 nsew signal output
rlabel metal2 s 8036 100 8148 400 6 la_data_out[2]
port 117 nsew signal output
rlabel metal2 s 8036 29600 8148 29900 6 la_data_out[30]
port 118 nsew signal output
rlabel metal3 s 29600 15092 29900 15204 6 la_data_out[31]
port 119 nsew signal output
rlabel metal2 s 4676 29600 4788 29900 6 la_data_out[32]
port 120 nsew signal output
rlabel metal3 s 29600 20132 29900 20244 6 la_data_out[33]
port 121 nsew signal output
rlabel metal3 s 100 29204 400 29316 6 la_data_out[34]
port 122 nsew signal output
rlabel metal3 s 100 23492 400 23604 6 la_data_out[35]
port 123 nsew signal output
rlabel metal3 s 29600 23156 29900 23268 6 la_data_out[36]
port 124 nsew signal output
rlabel metal3 s 29600 25508 29900 25620 6 la_data_out[37]
port 125 nsew signal output
rlabel metal3 s 100 9716 400 9828 6 la_data_out[38]
port 126 nsew signal output
rlabel metal2 s 25508 100 25620 400 6 la_data_out[39]
port 127 nsew signal output
rlabel metal3 s 100 15428 400 15540 6 la_data_out[3]
port 128 nsew signal output
rlabel metal3 s 29600 29204 29900 29316 6 la_data_out[40]
port 129 nsew signal output
rlabel metal3 s 100 25508 400 25620 6 la_data_out[41]
port 130 nsew signal output
rlabel metal3 s 29600 12068 29900 12180 6 la_data_out[42]
port 131 nsew signal output
rlabel metal3 s 100 26852 400 26964 6 la_data_out[43]
port 132 nsew signal output
rlabel metal2 s 9380 100 9492 400 6 la_data_out[44]
port 133 nsew signal output
rlabel metal3 s 100 2324 400 2436 6 la_data_out[45]
port 134 nsew signal output
rlabel metal3 s 29600 19460 29900 19572 6 la_data_out[46]
port 135 nsew signal output
rlabel metal2 s 6692 29600 6804 29900 6 la_data_out[47]
port 136 nsew signal output
rlabel metal2 s 29876 29600 29988 29900 6 la_data_out[48]
port 137 nsew signal output
rlabel metal3 s 100 9044 400 9156 6 la_data_out[49]
port 138 nsew signal output
rlabel metal3 s 29600 5348 29900 5460 6 la_data_out[4]
port 139 nsew signal output
rlabel metal2 s 15764 29600 15876 29900 6 la_data_out[50]
port 140 nsew signal output
rlabel metal2 s 1652 100 1764 400 6 la_data_out[51]
port 141 nsew signal output
rlabel metal2 s 25172 100 25284 400 6 la_data_out[52]
port 142 nsew signal output
rlabel metal3 s 100 22484 400 22596 6 la_data_out[53]
port 143 nsew signal output
rlabel metal3 s 100 28532 400 28644 6 la_data_out[54]
port 144 nsew signal output
rlabel metal2 s 12068 100 12180 400 6 la_data_out[55]
port 145 nsew signal output
rlabel metal2 s 20468 29600 20580 29900 6 la_data_out[56]
port 146 nsew signal output
rlabel metal3 s 29600 23828 29900 23940 6 la_data_out[57]
port 147 nsew signal output
rlabel metal2 s 6356 29600 6468 29900 6 la_data_out[58]
port 148 nsew signal output
rlabel metal3 s 29600 15428 29900 15540 6 la_data_out[59]
port 149 nsew signal output
rlabel metal3 s 100 19460 400 19572 6 la_data_out[5]
port 150 nsew signal output
rlabel metal3 s 100 5012 400 5124 6 la_data_out[60]
port 151 nsew signal output
rlabel metal3 s 100 4676 400 4788 6 la_data_out[61]
port 152 nsew signal output
rlabel metal2 s 18452 29600 18564 29900 6 la_data_out[62]
port 153 nsew signal output
rlabel metal2 s 10388 29600 10500 29900 6 la_data_out[63]
port 154 nsew signal output
rlabel metal3 s 29600 980 29900 1092 6 la_data_out[6]
port 155 nsew signal output
rlabel metal2 s 13412 29600 13524 29900 6 la_data_out[7]
port 156 nsew signal output
rlabel metal2 s 5684 29600 5796 29900 6 la_data_out[8]
port 157 nsew signal output
rlabel metal3 s 100 26180 400 26292 6 la_data_out[9]
port 158 nsew signal output
rlabel metal3 s 29600 3668 29900 3780 6 la_oenb[0]
port 159 nsew signal input
rlabel metal3 s 100 15092 400 15204 6 la_oenb[10]
port 160 nsew signal input
rlabel metal3 s 29600 8708 29900 8820 6 la_oenb[11]
port 161 nsew signal input
rlabel metal2 s 18788 100 18900 400 6 la_oenb[12]
port 162 nsew signal input
rlabel metal2 s 17444 29600 17556 29900 6 la_oenb[13]
port 163 nsew signal input
rlabel metal2 s 18452 100 18564 400 6 la_oenb[14]
port 164 nsew signal input
rlabel metal3 s 100 644 400 756 6 la_oenb[15]
port 165 nsew signal input
rlabel metal2 s 3332 100 3444 400 6 la_oenb[16]
port 166 nsew signal input
rlabel metal2 s 5348 100 5460 400 6 la_oenb[17]
port 167 nsew signal input
rlabel metal2 s 22148 29600 22260 29900 6 la_oenb[18]
port 168 nsew signal input
rlabel metal2 s 21140 29600 21252 29900 6 la_oenb[19]
port 169 nsew signal input
rlabel metal3 s 100 5684 400 5796 6 la_oenb[1]
port 170 nsew signal input
rlabel metal3 s 29600 22484 29900 22596 6 la_oenb[20]
port 171 nsew signal input
rlabel metal3 s 100 2660 400 2772 6 la_oenb[21]
port 172 nsew signal input
rlabel metal3 s 100 18452 400 18564 6 la_oenb[22]
port 173 nsew signal input
rlabel metal2 s 7028 100 7140 400 6 la_oenb[23]
port 174 nsew signal input
rlabel metal2 s 11732 29600 11844 29900 6 la_oenb[24]
port 175 nsew signal input
rlabel metal2 s 1988 29600 2100 29900 6 la_oenb[25]
port 176 nsew signal input
rlabel metal3 s 100 5348 400 5460 6 la_oenb[26]
port 177 nsew signal input
rlabel metal3 s 100 9380 400 9492 6 la_oenb[27]
port 178 nsew signal input
rlabel metal3 s 29600 9044 29900 9156 6 la_oenb[28]
port 179 nsew signal input
rlabel metal3 s 29600 19796 29900 19908 6 la_oenb[29]
port 180 nsew signal input
rlabel metal3 s 29600 21812 29900 21924 6 la_oenb[2]
port 181 nsew signal input
rlabel metal3 s 29600 17780 29900 17892 6 la_oenb[30]
port 182 nsew signal input
rlabel metal2 s 23828 29600 23940 29900 6 la_oenb[31]
port 183 nsew signal input
rlabel metal3 s 29600 16772 29900 16884 6 la_oenb[32]
port 184 nsew signal input
rlabel metal2 s 13076 100 13188 400 6 la_oenb[33]
port 185 nsew signal input
rlabel metal3 s 29600 24500 29900 24612 6 la_oenb[34]
port 186 nsew signal input
rlabel metal3 s 100 13076 400 13188 6 la_oenb[35]
port 187 nsew signal input
rlabel metal2 s 308 100 420 400 6 la_oenb[36]
port 188 nsew signal input
rlabel metal2 s 17780 29600 17892 29900 6 la_oenb[37]
port 189 nsew signal input
rlabel metal2 s 13412 100 13524 400 6 la_oenb[38]
port 190 nsew signal input
rlabel metal2 s 27188 100 27300 400 6 la_oenb[39]
port 191 nsew signal input
rlabel metal3 s 100 25172 400 25284 6 la_oenb[3]
port 192 nsew signal input
rlabel metal2 s 29204 100 29316 400 6 la_oenb[40]
port 193 nsew signal input
rlabel metal2 s 20804 29600 20916 29900 6 la_oenb[41]
port 194 nsew signal input
rlabel metal3 s 100 23828 400 23940 6 la_oenb[42]
port 195 nsew signal input
rlabel metal2 s 5012 100 5124 400 6 la_oenb[43]
port 196 nsew signal input
rlabel metal3 s 100 4340 400 4452 6 la_oenb[44]
port 197 nsew signal input
rlabel metal3 s 29600 27188 29900 27300 6 la_oenb[45]
port 198 nsew signal input
rlabel metal2 s 20804 100 20916 400 6 la_oenb[46]
port 199 nsew signal input
rlabel metal2 s 10052 100 10164 400 6 la_oenb[47]
port 200 nsew signal input
rlabel metal3 s 100 16436 400 16548 6 la_oenb[48]
port 201 nsew signal input
rlabel metal3 s 29600 9380 29900 9492 6 la_oenb[49]
port 202 nsew signal input
rlabel metal2 s 4340 29600 4452 29900 6 la_oenb[4]
port 203 nsew signal input
rlabel metal2 s 20468 100 20580 400 6 la_oenb[50]
port 204 nsew signal input
rlabel metal2 s 18788 29600 18900 29900 6 la_oenb[51]
port 205 nsew signal input
rlabel metal2 s 26516 100 26628 400 6 la_oenb[52]
port 206 nsew signal input
rlabel metal3 s 100 23156 400 23268 6 la_oenb[53]
port 207 nsew signal input
rlabel metal3 s 100 24164 400 24276 6 la_oenb[54]
port 208 nsew signal input
rlabel metal3 s 29600 10388 29900 10500 6 la_oenb[55]
port 209 nsew signal input
rlabel metal2 s 20132 100 20244 400 6 la_oenb[56]
port 210 nsew signal input
rlabel metal3 s 29600 26852 29900 26964 6 la_oenb[57]
port 211 nsew signal input
rlabel metal2 s 29540 100 29652 400 6 la_oenb[58]
port 212 nsew signal input
rlabel metal2 s 25172 29600 25284 29900 6 la_oenb[59]
port 213 nsew signal input
rlabel metal2 s 24836 100 24948 400 6 la_oenb[5]
port 214 nsew signal input
rlabel metal2 s 15428 29600 15540 29900 6 la_oenb[60]
port 215 nsew signal input
rlabel metal2 s 2996 100 3108 400 6 la_oenb[61]
port 216 nsew signal input
rlabel metal3 s 29600 10724 29900 10836 6 la_oenb[62]
port 217 nsew signal input
rlabel metal2 s 980 29600 1092 29900 6 la_oenb[63]
port 218 nsew signal input
rlabel metal3 s 100 308 400 420 6 la_oenb[6]
port 219 nsew signal input
rlabel metal2 s 6692 100 6804 400 6 la_oenb[7]
port 220 nsew signal input
rlabel metal2 s 26180 100 26292 400 6 la_oenb[8]
port 221 nsew signal input
rlabel metal2 s 16100 29600 16212 29900 6 la_oenb[9]
port 222 nsew signal input
rlabel metal3 s 29600 28532 29900 28644 6 user_clock2
port 223 nsew signal input
rlabel metal3 s 100 20132 400 20244 6 user_irq[0]
port 224 nsew signal output
rlabel metal2 s 14756 29600 14868 29900 6 user_irq[1]
port 225 nsew signal output
rlabel metal2 s 16772 29600 16884 29900 6 user_irq[2]
port 226 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 227 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 227 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 228 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 228 nsew ground bidirectional
rlabel metal3 s 29600 1988 29900 2100 6 wb_clk_i
port 229 nsew signal input
rlabel metal2 s 12404 29600 12516 29900 6 wb_rst_i
port 230 nsew signal input
rlabel metal3 s 29600 6692 29900 6804 6 wbs_ack_o
port 231 nsew signal output
rlabel metal3 s 100 14756 400 14868 6 wbs_adr_i[0]
port 232 nsew signal input
rlabel metal2 s 19796 29600 19908 29900 6 wbs_adr_i[10]
port 233 nsew signal input
rlabel metal2 s 9044 29600 9156 29900 6 wbs_adr_i[11]
port 234 nsew signal input
rlabel metal2 s 2324 100 2436 400 6 wbs_adr_i[12]
port 235 nsew signal input
rlabel metal2 s 15428 100 15540 400 6 wbs_adr_i[13]
port 236 nsew signal input
rlabel metal3 s 29600 18116 29900 18228 6 wbs_adr_i[14]
port 237 nsew signal input
rlabel metal3 s 100 17780 400 17892 6 wbs_adr_i[15]
port 238 nsew signal input
rlabel metal2 s 17780 100 17892 400 6 wbs_adr_i[16]
port 239 nsew signal input
rlabel metal3 s 100 24500 400 24612 6 wbs_adr_i[17]
port 240 nsew signal input
rlabel metal3 s 29600 6356 29900 6468 6 wbs_adr_i[18]
port 241 nsew signal input
rlabel metal2 s 26852 100 26964 400 6 wbs_adr_i[19]
port 242 nsew signal input
rlabel metal3 s 100 12068 400 12180 6 wbs_adr_i[1]
port 243 nsew signal input
rlabel metal3 s 29600 27860 29900 27972 6 wbs_adr_i[20]
port 244 nsew signal input
rlabel metal2 s 15764 100 15876 400 6 wbs_adr_i[21]
port 245 nsew signal input
rlabel metal2 s 22820 100 22932 400 6 wbs_adr_i[22]
port 246 nsew signal input
rlabel metal3 s 29600 4340 29900 4452 6 wbs_adr_i[23]
port 247 nsew signal input
rlabel metal3 s 100 8708 400 8820 6 wbs_adr_i[24]
port 248 nsew signal input
rlabel metal2 s 15092 100 15204 400 6 wbs_adr_i[25]
port 249 nsew signal input
rlabel metal2 s 2660 100 2772 400 6 wbs_adr_i[26]
port 250 nsew signal input
rlabel metal2 s 15092 29600 15204 29900 6 wbs_adr_i[27]
port 251 nsew signal input
rlabel metal3 s 29600 14420 29900 14532 6 wbs_adr_i[28]
port 252 nsew signal input
rlabel metal3 s 100 14420 400 14532 6 wbs_adr_i[29]
port 253 nsew signal input
rlabel metal2 s 10724 100 10836 400 6 wbs_adr_i[2]
port 254 nsew signal input
rlabel metal2 s 27860 29600 27972 29900 6 wbs_adr_i[30]
port 255 nsew signal input
rlabel metal3 s 29600 10052 29900 10164 6 wbs_adr_i[31]
port 256 nsew signal input
rlabel metal2 s 22148 100 22260 400 6 wbs_adr_i[3]
port 257 nsew signal input
rlabel metal2 s 26852 29600 26964 29900 6 wbs_adr_i[4]
port 258 nsew signal input
rlabel metal2 s 21140 100 21252 400 6 wbs_adr_i[5]
port 259 nsew signal input
rlabel metal3 s 100 18116 400 18228 6 wbs_adr_i[6]
port 260 nsew signal input
rlabel metal2 s 1316 100 1428 400 6 wbs_adr_i[7]
port 261 nsew signal input
rlabel metal2 s 28532 100 28644 400 6 wbs_adr_i[8]
port 262 nsew signal input
rlabel metal3 s 29600 6020 29900 6132 6 wbs_adr_i[9]
port 263 nsew signal input
rlabel metal2 s 13748 29600 13860 29900 6 wbs_cyc_i
port 264 nsew signal input
rlabel metal3 s 29600 23492 29900 23604 6 wbs_dat_i[0]
port 265 nsew signal input
rlabel metal3 s 100 1988 400 2100 6 wbs_dat_i[10]
port 266 nsew signal input
rlabel metal3 s 100 29876 400 29988 6 wbs_dat_i[11]
port 267 nsew signal input
rlabel metal3 s 100 28868 400 28980 6 wbs_dat_i[12]
port 268 nsew signal input
rlabel metal2 s 980 100 1092 400 6 wbs_dat_i[13]
port 269 nsew signal input
rlabel metal3 s 100 7700 400 7812 6 wbs_dat_i[14]
port 270 nsew signal input
rlabel metal3 s 29600 13748 29900 13860 6 wbs_dat_i[15]
port 271 nsew signal input
rlabel metal2 s 16436 100 16548 400 6 wbs_dat_i[16]
port 272 nsew signal input
rlabel metal2 s 23492 29600 23604 29900 6 wbs_dat_i[17]
port 273 nsew signal input
rlabel metal3 s 29600 29540 29900 29652 6 wbs_dat_i[18]
port 274 nsew signal input
rlabel metal2 s 5348 29600 5460 29900 6 wbs_dat_i[19]
port 275 nsew signal input
rlabel metal2 s 4340 100 4452 400 6 wbs_dat_i[1]
port 276 nsew signal input
rlabel metal3 s 29600 16100 29900 16212 6 wbs_dat_i[20]
port 277 nsew signal input
rlabel metal3 s 29600 28868 29900 28980 6 wbs_dat_i[21]
port 278 nsew signal input
rlabel metal3 s 100 21812 400 21924 6 wbs_dat_i[22]
port 279 nsew signal input
rlabel metal3 s 29600 21140 29900 21252 6 wbs_dat_i[23]
port 280 nsew signal input
rlabel metal3 s 29600 8036 29900 8148 6 wbs_dat_i[24]
port 281 nsew signal input
rlabel metal3 s 100 11060 400 11172 6 wbs_dat_i[25]
port 282 nsew signal input
rlabel metal2 s 27524 29600 27636 29900 6 wbs_dat_i[26]
port 283 nsew signal input
rlabel metal2 s 10052 29600 10164 29900 6 wbs_dat_i[27]
port 284 nsew signal input
rlabel metal2 s 9044 100 9156 400 6 wbs_dat_i[28]
port 285 nsew signal input
rlabel metal3 s 29600 16436 29900 16548 6 wbs_dat_i[29]
port 286 nsew signal input
rlabel metal2 s 23828 100 23940 400 6 wbs_dat_i[2]
port 287 nsew signal input
rlabel metal3 s 29600 7364 29900 7476 6 wbs_dat_i[30]
port 288 nsew signal input
rlabel metal3 s 100 19124 400 19236 6 wbs_dat_i[31]
port 289 nsew signal input
rlabel metal3 s 29600 308 29900 420 6 wbs_dat_i[3]
port 290 nsew signal input
rlabel metal2 s 4676 100 4788 400 6 wbs_dat_i[4]
port 291 nsew signal input
rlabel metal2 s 14420 100 14532 400 6 wbs_dat_i[5]
port 292 nsew signal input
rlabel metal3 s 29600 11732 29900 11844 6 wbs_dat_i[6]
port 293 nsew signal input
rlabel metal2 s 25508 29600 25620 29900 6 wbs_dat_i[7]
port 294 nsew signal input
rlabel metal3 s 29600 25172 29900 25284 6 wbs_dat_i[8]
port 295 nsew signal input
rlabel metal3 s 29600 644 29900 756 6 wbs_dat_i[9]
port 296 nsew signal input
rlabel metal3 s 100 7364 400 7476 6 wbs_dat_o[0]
port 297 nsew signal output
rlabel metal3 s 29600 15764 29900 15876 6 wbs_dat_o[10]
port 298 nsew signal output
rlabel metal2 s 644 100 756 400 6 wbs_dat_o[11]
port 299 nsew signal output
rlabel metal3 s 29600 26516 29900 26628 6 wbs_dat_o[12]
port 300 nsew signal output
rlabel metal2 s 24164 29600 24276 29900 6 wbs_dat_o[13]
port 301 nsew signal output
rlabel metal3 s 29600 2660 29900 2772 6 wbs_dat_o[14]
port 302 nsew signal output
rlabel metal2 s 23156 29600 23268 29900 6 wbs_dat_o[15]
port 303 nsew signal output
rlabel metal3 s 100 10388 400 10500 6 wbs_dat_o[16]
port 304 nsew signal output
rlabel metal3 s 100 8036 400 8148 6 wbs_dat_o[17]
port 305 nsew signal output
rlabel metal2 s 19796 100 19908 400 6 wbs_dat_o[18]
port 306 nsew signal output
rlabel metal2 s -28 100 84 400 6 wbs_dat_o[19]
port 307 nsew signal output
rlabel metal2 s 23156 100 23268 400 6 wbs_dat_o[1]
port 308 nsew signal output
rlabel metal3 s 100 15764 400 15876 6 wbs_dat_o[20]
port 309 nsew signal output
rlabel metal3 s 100 27524 400 27636 6 wbs_dat_o[21]
port 310 nsew signal output
rlabel metal2 s 9380 29600 9492 29900 6 wbs_dat_o[22]
port 311 nsew signal output
rlabel metal3 s 100 11396 400 11508 6 wbs_dat_o[23]
port 312 nsew signal output
rlabel metal2 s 6020 100 6132 400 6 wbs_dat_o[24]
port 313 nsew signal output
rlabel metal2 s 1988 100 2100 400 6 wbs_dat_o[25]
port 314 nsew signal output
rlabel metal2 s 16436 29600 16548 29900 6 wbs_dat_o[26]
port 315 nsew signal output
rlabel metal2 s 9716 29600 9828 29900 6 wbs_dat_o[27]
port 316 nsew signal output
rlabel metal2 s 16100 100 16212 400 6 wbs_dat_o[28]
port 317 nsew signal output
rlabel metal2 s 21812 29600 21924 29900 6 wbs_dat_o[29]
port 318 nsew signal output
rlabel metal3 s 29600 7700 29900 7812 6 wbs_dat_o[2]
port 319 nsew signal output
rlabel metal3 s 100 20468 400 20580 6 wbs_dat_o[30]
port 320 nsew signal output
rlabel metal3 s 29600 22820 29900 22932 6 wbs_dat_o[31]
port 321 nsew signal output
rlabel metal2 s 6356 100 6468 400 6 wbs_dat_o[3]
port 322 nsew signal output
rlabel metal2 s 11396 100 11508 400 6 wbs_dat_o[4]
port 323 nsew signal output
rlabel metal3 s 100 2996 400 3108 6 wbs_dat_o[5]
port 324 nsew signal output
rlabel metal3 s 29600 22148 29900 22260 6 wbs_dat_o[6]
port 325 nsew signal output
rlabel metal2 s 18116 100 18228 400 6 wbs_dat_o[7]
port 326 nsew signal output
rlabel metal2 s 20132 29600 20244 29900 6 wbs_dat_o[8]
port 327 nsew signal output
rlabel metal2 s 19460 29600 19572 29900 6 wbs_dat_o[9]
port 328 nsew signal output
rlabel metal3 s 100 28196 400 28308 6 wbs_sel_i[0]
port 329 nsew signal input
rlabel metal2 s 2996 29600 3108 29900 6 wbs_sel_i[1]
port 330 nsew signal input
rlabel metal2 s 21812 100 21924 400 6 wbs_sel_i[2]
port 331 nsew signal input
rlabel metal3 s 100 6692 400 6804 6 wbs_sel_i[3]
port 332 nsew signal input
rlabel metal3 s 100 24836 400 24948 6 wbs_stb_i
port 333 nsew signal input
rlabel metal3 s 29600 14756 29900 14868 6 wbs_we_i
port 334 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 833780
string GDS_FILE /root/gf180-demo/caravel_user_project/openlane/top_wrapper/runs/22_12_03_21_00/results/signoff/top_wrapper.magic.gds
string GDS_START 156436
<< end >>

