VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_wrapper
  CLASS BLOCK ;
  FOREIGN top_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 184.520 299.000 185.640 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 241.640 299.000 242.760 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 296.000 27.720 299.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.040 296.000 293.160 299.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.840 1.000 141.960 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 113.960 299.000 115.080 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.200 296.000 229.320 299.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.400 296.000 296.520 299.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 97.160 299.000 98.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.840 1.000 57.960 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 261.800 299.000 262.920 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.600 296.000 111.720 299.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 9.800 4.000 10.920 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 70.280 4.000 71.400 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 197.960 4.000 199.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.600 1.000 195.720 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.240 296.000 24.360 299.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.160 296.000 182.280 299.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.440 1.000 175.560 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 63.560 4.000 64.680 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 265.160 4.000 266.280 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 204.680 299.000 205.800 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 271.880 4.000 273.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.000 1.000 246.120 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 248.360 299.000 249.480 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.040 4.000 125.160 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.160 296.000 14.280 299.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 174.440 299.000 175.560 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.960 296.000 283.080 299.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.200 296.000 61.320 299.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 134.120 299.000 135.240 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.880 1.000 105.000 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 23.240 299.000 24.360 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 110.600 299.000 111.720 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.320 296.000 286.440 299.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.560 1.000 148.680 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 124.040 299.000 125.160 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.080 296.000 4.200 299.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 295.400 4.000 296.520 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.080 1.000 88.200 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.840 1.000 225.960 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.840 296.000 225.960 299.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 296.000 115.080 299.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 130.760 299.000 131.880 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 137.480 4.000 138.600 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.120 296.000 51.240 299.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.320 1.000 118.440 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 296.000 145.320 299.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 208.040 299.000 209.160 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.160 296.000 266.280 299.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 117.320 4.000 118.440 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 33.320 299.000 34.440 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 278.600 4.000 279.720 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 281.960 299.000 283.080 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 187.880 299.000 189.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.040 4.000 209.160 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.240 1.000 276.360 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 46.760 299.000 47.880 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.360 296.000 249.480 299.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.680 296.000 37.800 299.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.800 296.000 262.920 299.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 187.880 4.000 189.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.640 296.000 74.760 299.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 13.160 4.000 14.280 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.760 296.000 131.880 299.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.000 1.000 78.120 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 50.120 299.000 51.240 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.880 296.000 273.000 299.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.720 1.000 168.840 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 191.240 299.000 192.360 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.320 4.000 34.440 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 29.960 299.000 31.080 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.480 1.000 138.600 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.200 4.000 61.320 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 211.400 4.000 212.520 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 16.520 4.000 17.640 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 161.000 4.000 162.120 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.080 296.000 88.200 299.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 13.160 299.000 14.280 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 70.280 299.000 71.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 100.520 4.000 101.640 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.040 1.000 125.160 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.240 1.000 192.360 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.240 296.000 108.360 299.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 275.240 299.000 276.360 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.680 296.000 121.800 299.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.960 1.000 283.080 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.160 1.000 98.280 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 167.720 4.000 168.840 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 56.840 299.000 57.960 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.680 1.000 37.800 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.320 296.000 34.440 299.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.000 296.000 78.120 299.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 36.680 4.000 37.800 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 -0.280 299.000 0.840 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 296.000 289.800 299.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.120 4.000 135.240 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.240 4.000 108.360 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.640 1.000 74.760 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.680 1.000 289.800 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.200 4.000 229.320 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 16.520 299.000 17.640 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.480 4.000 222.600 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.920 1.000 236.040 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.600 1.000 111.720 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 140.840 4.000 141.960 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 174.440 4.000 175.560 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.840 296.000 141.960 299.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.520 296.000 17.640 299.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 140.840 299.000 141.960 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.600 1.000 279.720 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.240 296.000 192.360 299.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.640 1.000 242.760 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.440 296.000 7.560 299.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.280 296.000 71.400 299.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.000 296.000 246.120 299.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 1.000 81.480 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.360 296.000 81.480 299.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 150.920 299.000 152.040 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.760 296.000 47.880 299.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 201.320 299.000 202.440 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 292.040 4.000 293.160 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 234.920 4.000 236.040 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 231.560 299.000 232.680 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 255.080 299.000 256.200 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 97.160 4.000 98.280 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.080 1.000 256.200 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 154.280 4.000 155.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 292.040 299.000 293.160 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 255.080 4.000 256.200 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 120.680 299.000 121.800 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 268.520 4.000 269.640 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.800 1.000 94.920 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 23.240 4.000 24.360 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 194.600 299.000 195.720 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.920 296.000 68.040 299.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 298.760 296.000 299.880 299.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 90.440 4.000 91.560 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 53.480 299.000 54.600 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.640 296.000 158.760 299.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.520 1.000 17.640 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.720 1.000 252.840 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 224.840 4.000 225.960 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 285.320 4.000 286.440 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.680 1.000 121.800 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.680 296.000 205.800 299.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 238.280 299.000 239.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.560 296.000 64.680 299.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 154.280 299.000 155.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.600 4.000 195.720 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 50.120 4.000 51.240 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 46.760 4.000 47.880 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.520 296.000 185.640 299.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.880 296.000 105.000 299.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 9.800 299.000 10.920 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.120 296.000 135.240 299.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.840 296.000 57.960 299.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 261.800 4.000 262.920 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 36.680 299.000 37.800 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 150.920 4.000 152.040 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 87.080 299.000 88.200 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.880 1.000 189.000 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.440 296.000 175.560 299.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.520 1.000 185.640 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 6.440 4.000 7.560 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.320 1.000 34.440 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 1.000 54.600 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.480 296.000 222.600 299.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.400 296.000 212.520 299.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 56.840 4.000 57.960 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 224.840 299.000 225.960 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.600 4.000 27.720 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 184.520 4.000 185.640 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.280 1.000 71.400 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.320 296.000 118.440 299.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.880 296.000 21.000 299.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.480 4.000 54.600 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 93.800 4.000 94.920 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 90.440 299.000 91.560 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 197.960 299.000 199.080 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 218.120 299.000 219.240 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 177.800 299.000 178.920 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.280 296.000 239.400 299.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 167.720 299.000 168.840 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 130.760 1.000 131.880 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 245.000 299.000 246.120 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 130.760 4.000 131.880 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.080 1.000 4.200 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.800 296.000 178.920 299.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.120 1.000 135.240 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.880 1.000 273.000 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 251.720 4.000 252.840 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.040 1.000 293.160 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.040 296.000 209.160 299.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 238.280 4.000 239.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.120 1.000 51.240 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 43.400 4.000 44.520 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 271.880 299.000 273.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.040 1.000 209.160 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.520 1.000 101.640 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 164.360 4.000 165.480 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 93.800 299.000 94.920 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.400 296.000 44.520 299.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.680 1.000 205.800 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.880 296.000 189.000 299.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 265.160 1.000 266.280 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 231.560 4.000 232.680 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 241.640 4.000 242.760 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 103.880 299.000 105.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.320 1.000 202.440 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 268.520 299.000 269.640 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.400 1.000 296.520 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 251.720 296.000 252.840 299.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.360 1.000 249.480 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.280 296.000 155.400 299.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.960 1.000 31.080 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 107.240 299.000 108.360 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.800 296.000 10.920 299.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 3.080 4.000 4.200 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.920 1.000 68.040 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 261.800 1.000 262.920 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.000 296.000 162.120 299.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 285.320 299.000 286.440 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 201.320 4.000 202.440 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.560 296.000 148.680 299.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 167.720 296.000 168.840 299.000 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 19.880 299.000 21.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.040 296.000 125.160 299.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 66.920 299.000 68.040 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 147.560 4.000 148.680 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.960 296.000 199.080 299.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.440 296.000 91.560 299.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.240 1.000 24.360 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.280 1.000 155.400 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 181.160 299.000 182.280 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 177.800 4.000 178.920 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 177.800 1.000 178.920 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 245.000 4.000 246.120 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 63.560 299.000 64.680 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.520 1.000 269.640 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 120.680 4.000 121.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 278.600 299.000 279.720 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.640 1.000 158.760 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.200 1.000 229.320 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 43.400 299.000 44.520 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 87.080 4.000 88.200 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.920 1.000 152.040 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.600 1.000 27.720 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.920 296.000 152.040 299.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 144.200 299.000 145.320 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.200 4.000 145.320 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.240 1.000 108.360 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.600 296.000 279.720 299.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 100.520 299.000 101.640 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.480 1.000 222.600 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.520 296.000 269.640 299.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.400 1.000 212.520 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 181.160 4.000 182.280 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.160 1.000 14.280 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.320 1.000 286.440 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 60.200 299.000 61.320 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.480 296.000 138.600 299.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 234.920 299.000 236.040 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 19.880 4.000 21.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 298.760 4.000 299.880 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.680 4.000 289.800 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 9.800 1.000 10.920 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 77.000 4.000 78.120 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 137.480 299.000 138.600 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.360 1.000 165.480 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.920 296.000 236.040 299.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 295.400 299.000 296.520 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.480 296.000 54.600 299.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.400 1.000 44.520 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 161.000 299.000 162.120 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 288.680 299.000 289.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.120 4.000 219.240 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 211.400 299.000 212.520 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 80.360 299.000 81.480 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 110.600 4.000 111.720 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.240 296.000 276.360 299.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.520 296.000 101.640 299.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.440 1.000 91.560 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 164.360 299.000 165.480 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.280 1.000 239.400 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 73.640 299.000 74.760 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.240 4.000 192.360 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 3.080 299.000 4.200 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 46.760 1.000 47.880 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.200 1.000 145.320 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 117.320 299.000 118.440 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.080 296.000 256.200 299.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 251.720 299.000 252.840 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 6.440 299.000 7.560 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 73.640 4.000 74.760 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 157.640 299.000 158.760 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.440 1.000 7.560 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 265.160 299.000 266.280 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.640 296.000 242.760 299.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 26.600 299.000 27.720 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.560 296.000 232.680 299.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 103.880 4.000 105.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 80.360 4.000 81.480 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.960 1.000 199.080 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT -0.280 1.000 0.840 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.560 1.000 232.680 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 157.640 4.000 158.760 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.240 4.000 276.360 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 93.800 296.000 94.920 299.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 113.960 4.000 115.080 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.200 1.000 61.320 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.880 1.000 21.000 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.360 296.000 165.480 299.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.160 296.000 98.280 299.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.000 1.000 162.120 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 296.000 219.240 299.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 77.000 299.000 78.120 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 204.680 4.000 205.800 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 228.200 299.000 229.320 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 63.560 1.000 64.680 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.960 1.000 115.080 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 29.960 4.000 31.080 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 221.480 299.000 222.600 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.160 1.000 182.280 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.320 296.000 202.440 299.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.600 296.000 195.720 299.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 281.960 4.000 283.080 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.960 296.000 31.080 299.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.120 1.000 219.240 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 66.920 4.000 68.040 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.360 4.000 249.480 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 147.560 299.000 148.680 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 292.880 283.770 ;
      LAYER Metal2 ;
        RECT 0.700 295.700 2.780 296.660 ;
        RECT 4.500 295.700 6.140 296.660 ;
        RECT 7.860 295.700 9.500 296.660 ;
        RECT 11.220 295.700 12.860 296.660 ;
        RECT 14.580 295.700 16.220 296.660 ;
        RECT 17.940 295.700 19.580 296.660 ;
        RECT 21.300 295.700 22.940 296.660 ;
        RECT 24.660 295.700 26.300 296.660 ;
        RECT 28.020 295.700 29.660 296.660 ;
        RECT 31.380 295.700 33.020 296.660 ;
        RECT 34.740 295.700 36.380 296.660 ;
        RECT 38.100 295.700 43.100 296.660 ;
        RECT 44.820 295.700 46.460 296.660 ;
        RECT 48.180 295.700 49.820 296.660 ;
        RECT 51.540 295.700 53.180 296.660 ;
        RECT 54.900 295.700 56.540 296.660 ;
        RECT 58.260 295.700 59.900 296.660 ;
        RECT 61.620 295.700 63.260 296.660 ;
        RECT 64.980 295.700 66.620 296.660 ;
        RECT 68.340 295.700 69.980 296.660 ;
        RECT 71.700 295.700 73.340 296.660 ;
        RECT 75.060 295.700 76.700 296.660 ;
        RECT 78.420 295.700 80.060 296.660 ;
        RECT 81.780 295.700 86.780 296.660 ;
        RECT 88.500 295.700 90.140 296.660 ;
        RECT 91.860 295.700 93.500 296.660 ;
        RECT 95.220 295.700 96.860 296.660 ;
        RECT 98.580 295.700 100.220 296.660 ;
        RECT 101.940 295.700 103.580 296.660 ;
        RECT 105.300 295.700 106.940 296.660 ;
        RECT 108.660 295.700 110.300 296.660 ;
        RECT 112.020 295.700 113.660 296.660 ;
        RECT 115.380 295.700 117.020 296.660 ;
        RECT 118.740 295.700 120.380 296.660 ;
        RECT 122.100 295.700 123.740 296.660 ;
        RECT 125.460 295.700 130.460 296.660 ;
        RECT 132.180 295.700 133.820 296.660 ;
        RECT 135.540 295.700 137.180 296.660 ;
        RECT 138.900 295.700 140.540 296.660 ;
        RECT 142.260 295.700 143.900 296.660 ;
        RECT 145.620 295.700 147.260 296.660 ;
        RECT 148.980 295.700 150.620 296.660 ;
        RECT 152.340 295.700 153.980 296.660 ;
        RECT 155.700 295.700 157.340 296.660 ;
        RECT 159.060 295.700 160.700 296.660 ;
        RECT 162.420 295.700 164.060 296.660 ;
        RECT 165.780 295.700 167.420 296.660 ;
        RECT 169.140 295.700 174.140 296.660 ;
        RECT 175.860 295.700 177.500 296.660 ;
        RECT 179.220 295.700 180.860 296.660 ;
        RECT 182.580 295.700 184.220 296.660 ;
        RECT 185.940 295.700 187.580 296.660 ;
        RECT 189.300 295.700 190.940 296.660 ;
        RECT 192.660 295.700 194.300 296.660 ;
        RECT 196.020 295.700 197.660 296.660 ;
        RECT 199.380 295.700 201.020 296.660 ;
        RECT 202.740 295.700 204.380 296.660 ;
        RECT 206.100 295.700 207.740 296.660 ;
        RECT 209.460 295.700 211.100 296.660 ;
        RECT 212.820 295.700 217.820 296.660 ;
        RECT 219.540 295.700 221.180 296.660 ;
        RECT 222.900 295.700 224.540 296.660 ;
        RECT 226.260 295.700 227.900 296.660 ;
        RECT 229.620 295.700 231.260 296.660 ;
        RECT 232.980 295.700 234.620 296.660 ;
        RECT 236.340 295.700 237.980 296.660 ;
        RECT 239.700 295.700 241.340 296.660 ;
        RECT 243.060 295.700 244.700 296.660 ;
        RECT 246.420 295.700 248.060 296.660 ;
        RECT 249.780 295.700 251.420 296.660 ;
        RECT 253.140 295.700 254.780 296.660 ;
        RECT 256.500 295.700 261.500 296.660 ;
        RECT 263.220 295.700 264.860 296.660 ;
        RECT 266.580 295.700 268.220 296.660 ;
        RECT 269.940 295.700 271.580 296.660 ;
        RECT 273.300 295.700 274.940 296.660 ;
        RECT 276.660 295.700 278.300 296.660 ;
        RECT 280.020 295.700 281.660 296.660 ;
        RECT 283.380 295.700 285.020 296.660 ;
        RECT 286.740 295.700 288.380 296.660 ;
        RECT 290.100 295.700 291.740 296.660 ;
        RECT 293.460 295.700 295.100 296.660 ;
        RECT 296.820 295.700 298.460 296.660 ;
        RECT 0.700 4.300 298.900 295.700 ;
        RECT 1.140 0.700 2.780 4.300 ;
        RECT 4.500 0.700 6.140 4.300 ;
        RECT 7.860 0.700 9.500 4.300 ;
        RECT 11.220 0.700 12.860 4.300 ;
        RECT 14.580 0.700 16.220 4.300 ;
        RECT 17.940 0.700 19.580 4.300 ;
        RECT 21.300 0.700 22.940 4.300 ;
        RECT 24.660 0.700 26.300 4.300 ;
        RECT 28.020 0.700 29.660 4.300 ;
        RECT 31.380 0.700 33.020 4.300 ;
        RECT 34.740 0.700 36.380 4.300 ;
        RECT 38.100 0.700 43.100 4.300 ;
        RECT 44.820 0.700 46.460 4.300 ;
        RECT 48.180 0.700 49.820 4.300 ;
        RECT 51.540 0.700 53.180 4.300 ;
        RECT 54.900 0.700 56.540 4.300 ;
        RECT 58.260 0.700 59.900 4.300 ;
        RECT 61.620 0.700 63.260 4.300 ;
        RECT 64.980 0.700 66.620 4.300 ;
        RECT 68.340 0.700 69.980 4.300 ;
        RECT 71.700 0.700 73.340 4.300 ;
        RECT 75.060 0.700 76.700 4.300 ;
        RECT 78.420 0.700 80.060 4.300 ;
        RECT 81.780 0.700 86.780 4.300 ;
        RECT 88.500 0.700 90.140 4.300 ;
        RECT 91.860 0.700 93.500 4.300 ;
        RECT 95.220 0.700 96.860 4.300 ;
        RECT 98.580 0.700 100.220 4.300 ;
        RECT 101.940 0.700 103.580 4.300 ;
        RECT 105.300 0.700 106.940 4.300 ;
        RECT 108.660 0.700 110.300 4.300 ;
        RECT 112.020 0.700 113.660 4.300 ;
        RECT 115.380 0.700 117.020 4.300 ;
        RECT 118.740 0.700 120.380 4.300 ;
        RECT 122.100 0.700 123.740 4.300 ;
        RECT 125.460 0.700 130.460 4.300 ;
        RECT 132.180 0.700 133.820 4.300 ;
        RECT 135.540 0.700 137.180 4.300 ;
        RECT 138.900 0.700 140.540 4.300 ;
        RECT 142.260 0.700 143.900 4.300 ;
        RECT 145.620 0.700 147.260 4.300 ;
        RECT 148.980 0.700 150.620 4.300 ;
        RECT 152.340 0.700 153.980 4.300 ;
        RECT 155.700 0.700 157.340 4.300 ;
        RECT 159.060 0.700 160.700 4.300 ;
        RECT 162.420 0.700 164.060 4.300 ;
        RECT 165.780 0.700 167.420 4.300 ;
        RECT 169.140 0.700 174.140 4.300 ;
        RECT 175.860 0.700 177.500 4.300 ;
        RECT 179.220 0.700 180.860 4.300 ;
        RECT 182.580 0.700 184.220 4.300 ;
        RECT 185.940 0.700 187.580 4.300 ;
        RECT 189.300 0.700 190.940 4.300 ;
        RECT 192.660 0.700 194.300 4.300 ;
        RECT 196.020 0.700 197.660 4.300 ;
        RECT 199.380 0.700 201.020 4.300 ;
        RECT 202.740 0.700 204.380 4.300 ;
        RECT 206.100 0.700 207.740 4.300 ;
        RECT 209.460 0.700 211.100 4.300 ;
        RECT 212.820 0.700 217.820 4.300 ;
        RECT 219.540 0.700 221.180 4.300 ;
        RECT 222.900 0.700 224.540 4.300 ;
        RECT 226.260 0.700 227.900 4.300 ;
        RECT 229.620 0.700 231.260 4.300 ;
        RECT 232.980 0.700 234.620 4.300 ;
        RECT 236.340 0.700 237.980 4.300 ;
        RECT 239.700 0.700 241.340 4.300 ;
        RECT 243.060 0.700 244.700 4.300 ;
        RECT 246.420 0.700 248.060 4.300 ;
        RECT 249.780 0.700 251.420 4.300 ;
        RECT 253.140 0.700 254.780 4.300 ;
        RECT 256.500 0.700 261.500 4.300 ;
        RECT 263.220 0.700 264.860 4.300 ;
        RECT 266.580 0.700 268.220 4.300 ;
        RECT 269.940 0.700 271.580 4.300 ;
        RECT 273.300 0.700 274.940 4.300 ;
        RECT 276.660 0.700 278.300 4.300 ;
        RECT 280.020 0.700 281.660 4.300 ;
        RECT 283.380 0.700 285.020 4.300 ;
        RECT 286.740 0.700 288.380 4.300 ;
        RECT 290.100 0.700 291.740 4.300 ;
        RECT 293.460 0.700 295.100 4.300 ;
        RECT 296.820 0.700 298.900 4.300 ;
        RECT 0.700 0.650 298.900 0.700 ;
      LAYER Metal3 ;
        RECT 0.650 291.740 0.700 292.180 ;
        RECT 4.300 291.740 295.700 292.180 ;
        RECT 0.650 290.100 298.950 291.740 ;
        RECT 0.650 288.380 0.700 290.100 ;
        RECT 4.300 288.380 295.700 290.100 ;
        RECT 0.650 286.740 298.950 288.380 ;
        RECT 0.650 285.020 0.700 286.740 ;
        RECT 4.300 285.020 295.700 286.740 ;
        RECT 0.650 283.380 298.950 285.020 ;
        RECT 0.650 281.660 0.700 283.380 ;
        RECT 4.300 281.660 295.700 283.380 ;
        RECT 0.650 280.020 298.950 281.660 ;
        RECT 0.650 278.300 0.700 280.020 ;
        RECT 4.300 278.300 295.700 280.020 ;
        RECT 0.650 276.660 298.950 278.300 ;
        RECT 0.650 274.940 0.700 276.660 ;
        RECT 4.300 274.940 295.700 276.660 ;
        RECT 0.650 273.300 298.950 274.940 ;
        RECT 0.650 271.580 0.700 273.300 ;
        RECT 4.300 271.580 295.700 273.300 ;
        RECT 0.650 269.940 298.950 271.580 ;
        RECT 0.650 268.220 0.700 269.940 ;
        RECT 4.300 268.220 295.700 269.940 ;
        RECT 0.650 266.580 298.950 268.220 ;
        RECT 0.650 264.860 0.700 266.580 ;
        RECT 4.300 264.860 295.700 266.580 ;
        RECT 0.650 263.220 298.950 264.860 ;
        RECT 0.650 261.500 0.700 263.220 ;
        RECT 4.300 261.500 295.700 263.220 ;
        RECT 0.650 256.500 298.950 261.500 ;
        RECT 0.650 254.780 0.700 256.500 ;
        RECT 4.300 254.780 295.700 256.500 ;
        RECT 0.650 253.140 298.950 254.780 ;
        RECT 0.650 251.420 0.700 253.140 ;
        RECT 4.300 251.420 295.700 253.140 ;
        RECT 0.650 249.780 298.950 251.420 ;
        RECT 0.650 248.060 0.700 249.780 ;
        RECT 4.300 248.060 295.700 249.780 ;
        RECT 0.650 246.420 298.950 248.060 ;
        RECT 0.650 244.700 0.700 246.420 ;
        RECT 4.300 244.700 295.700 246.420 ;
        RECT 0.650 243.060 298.950 244.700 ;
        RECT 0.650 241.340 0.700 243.060 ;
        RECT 4.300 241.340 295.700 243.060 ;
        RECT 0.650 239.700 298.950 241.340 ;
        RECT 0.650 237.980 0.700 239.700 ;
        RECT 4.300 237.980 295.700 239.700 ;
        RECT 0.650 236.340 298.950 237.980 ;
        RECT 0.650 234.620 0.700 236.340 ;
        RECT 4.300 234.620 295.700 236.340 ;
        RECT 0.650 232.980 298.950 234.620 ;
        RECT 0.650 231.260 0.700 232.980 ;
        RECT 4.300 231.260 295.700 232.980 ;
        RECT 0.650 229.620 298.950 231.260 ;
        RECT 0.650 227.900 0.700 229.620 ;
        RECT 4.300 227.900 295.700 229.620 ;
        RECT 0.650 226.260 298.950 227.900 ;
        RECT 0.650 224.540 0.700 226.260 ;
        RECT 4.300 224.540 295.700 226.260 ;
        RECT 0.650 222.900 298.950 224.540 ;
        RECT 0.650 221.180 0.700 222.900 ;
        RECT 4.300 221.180 295.700 222.900 ;
        RECT 0.650 219.540 298.950 221.180 ;
        RECT 0.650 217.820 0.700 219.540 ;
        RECT 4.300 217.820 295.700 219.540 ;
        RECT 0.650 212.820 298.950 217.820 ;
        RECT 0.650 211.100 0.700 212.820 ;
        RECT 4.300 211.100 295.700 212.820 ;
        RECT 0.650 209.460 298.950 211.100 ;
        RECT 0.650 207.740 0.700 209.460 ;
        RECT 4.300 207.740 295.700 209.460 ;
        RECT 0.650 206.100 298.950 207.740 ;
        RECT 0.650 204.380 0.700 206.100 ;
        RECT 4.300 204.380 295.700 206.100 ;
        RECT 0.650 202.740 298.950 204.380 ;
        RECT 0.650 201.020 0.700 202.740 ;
        RECT 4.300 201.020 295.700 202.740 ;
        RECT 0.650 199.380 298.950 201.020 ;
        RECT 0.650 197.660 0.700 199.380 ;
        RECT 4.300 197.660 295.700 199.380 ;
        RECT 0.650 196.020 298.950 197.660 ;
        RECT 0.650 194.300 0.700 196.020 ;
        RECT 4.300 194.300 295.700 196.020 ;
        RECT 0.650 192.660 298.950 194.300 ;
        RECT 0.650 190.940 0.700 192.660 ;
        RECT 4.300 190.940 295.700 192.660 ;
        RECT 0.650 189.300 298.950 190.940 ;
        RECT 0.650 187.580 0.700 189.300 ;
        RECT 4.300 187.580 295.700 189.300 ;
        RECT 0.650 185.940 298.950 187.580 ;
        RECT 0.650 184.220 0.700 185.940 ;
        RECT 4.300 184.220 295.700 185.940 ;
        RECT 0.650 182.580 298.950 184.220 ;
        RECT 0.650 180.860 0.700 182.580 ;
        RECT 4.300 180.860 295.700 182.580 ;
        RECT 0.650 179.220 298.950 180.860 ;
        RECT 0.650 177.500 0.700 179.220 ;
        RECT 4.300 177.500 295.700 179.220 ;
        RECT 0.650 175.860 298.950 177.500 ;
        RECT 0.650 174.140 0.700 175.860 ;
        RECT 4.300 174.140 295.700 175.860 ;
        RECT 0.650 169.140 298.950 174.140 ;
        RECT 0.650 167.420 0.700 169.140 ;
        RECT 4.300 167.420 295.700 169.140 ;
        RECT 0.650 165.780 298.950 167.420 ;
        RECT 0.650 164.060 0.700 165.780 ;
        RECT 4.300 164.060 295.700 165.780 ;
        RECT 0.650 162.420 298.950 164.060 ;
        RECT 0.650 160.700 0.700 162.420 ;
        RECT 4.300 160.700 295.700 162.420 ;
        RECT 0.650 159.060 298.950 160.700 ;
        RECT 0.650 157.340 0.700 159.060 ;
        RECT 4.300 157.340 295.700 159.060 ;
        RECT 0.650 155.700 298.950 157.340 ;
        RECT 0.650 153.980 0.700 155.700 ;
        RECT 4.300 153.980 295.700 155.700 ;
        RECT 0.650 152.340 298.950 153.980 ;
        RECT 0.650 150.620 0.700 152.340 ;
        RECT 4.300 150.620 295.700 152.340 ;
        RECT 0.650 148.980 298.950 150.620 ;
        RECT 0.650 147.260 0.700 148.980 ;
        RECT 4.300 147.260 295.700 148.980 ;
        RECT 0.650 145.620 298.950 147.260 ;
        RECT 0.650 143.900 0.700 145.620 ;
        RECT 4.300 143.900 295.700 145.620 ;
        RECT 0.650 142.260 298.950 143.900 ;
        RECT 0.650 140.540 0.700 142.260 ;
        RECT 4.300 140.540 295.700 142.260 ;
        RECT 0.650 138.900 298.950 140.540 ;
        RECT 0.650 137.180 0.700 138.900 ;
        RECT 4.300 137.180 295.700 138.900 ;
        RECT 0.650 135.540 298.950 137.180 ;
        RECT 0.650 133.820 0.700 135.540 ;
        RECT 4.300 133.820 295.700 135.540 ;
        RECT 0.650 132.180 298.950 133.820 ;
        RECT 0.650 130.460 0.700 132.180 ;
        RECT 4.300 130.460 295.700 132.180 ;
        RECT 0.650 125.460 298.950 130.460 ;
        RECT 0.650 123.740 0.700 125.460 ;
        RECT 4.300 123.740 295.700 125.460 ;
        RECT 0.650 122.100 298.950 123.740 ;
        RECT 0.650 120.380 0.700 122.100 ;
        RECT 4.300 120.380 295.700 122.100 ;
        RECT 0.650 118.740 298.950 120.380 ;
        RECT 0.650 117.020 0.700 118.740 ;
        RECT 4.300 117.020 295.700 118.740 ;
        RECT 0.650 115.380 298.950 117.020 ;
        RECT 0.650 113.660 0.700 115.380 ;
        RECT 4.300 113.660 295.700 115.380 ;
        RECT 0.650 112.020 298.950 113.660 ;
        RECT 0.650 110.300 0.700 112.020 ;
        RECT 4.300 110.300 295.700 112.020 ;
        RECT 0.650 108.660 298.950 110.300 ;
        RECT 0.650 106.940 0.700 108.660 ;
        RECT 4.300 106.940 295.700 108.660 ;
        RECT 0.650 105.300 298.950 106.940 ;
        RECT 0.650 103.580 0.700 105.300 ;
        RECT 4.300 103.580 295.700 105.300 ;
        RECT 0.650 101.940 298.950 103.580 ;
        RECT 0.650 100.220 0.700 101.940 ;
        RECT 4.300 100.220 295.700 101.940 ;
        RECT 0.650 98.580 298.950 100.220 ;
        RECT 0.650 96.860 0.700 98.580 ;
        RECT 4.300 96.860 295.700 98.580 ;
        RECT 0.650 95.220 298.950 96.860 ;
        RECT 0.650 93.500 0.700 95.220 ;
        RECT 4.300 93.500 295.700 95.220 ;
        RECT 0.650 91.860 298.950 93.500 ;
        RECT 0.650 90.140 0.700 91.860 ;
        RECT 4.300 90.140 295.700 91.860 ;
        RECT 0.650 88.500 298.950 90.140 ;
        RECT 0.650 86.780 0.700 88.500 ;
        RECT 4.300 86.780 295.700 88.500 ;
        RECT 0.650 81.780 298.950 86.780 ;
        RECT 0.650 80.060 0.700 81.780 ;
        RECT 4.300 80.060 295.700 81.780 ;
        RECT 0.650 78.420 298.950 80.060 ;
        RECT 0.650 76.700 0.700 78.420 ;
        RECT 4.300 76.700 295.700 78.420 ;
        RECT 0.650 75.060 298.950 76.700 ;
        RECT 0.650 73.340 0.700 75.060 ;
        RECT 4.300 73.340 295.700 75.060 ;
        RECT 0.650 71.700 298.950 73.340 ;
        RECT 0.650 69.980 0.700 71.700 ;
        RECT 4.300 69.980 295.700 71.700 ;
        RECT 0.650 68.340 298.950 69.980 ;
        RECT 0.650 66.620 0.700 68.340 ;
        RECT 4.300 66.620 295.700 68.340 ;
        RECT 0.650 64.980 298.950 66.620 ;
        RECT 0.650 63.260 0.700 64.980 ;
        RECT 4.300 63.260 295.700 64.980 ;
        RECT 0.650 61.620 298.950 63.260 ;
        RECT 0.650 59.900 0.700 61.620 ;
        RECT 4.300 59.900 295.700 61.620 ;
        RECT 0.650 58.260 298.950 59.900 ;
        RECT 0.650 56.540 0.700 58.260 ;
        RECT 4.300 56.540 295.700 58.260 ;
        RECT 0.650 54.900 298.950 56.540 ;
        RECT 0.650 53.180 0.700 54.900 ;
        RECT 4.300 53.180 295.700 54.900 ;
        RECT 0.650 51.540 298.950 53.180 ;
        RECT 0.650 49.820 0.700 51.540 ;
        RECT 4.300 49.820 295.700 51.540 ;
        RECT 0.650 48.180 298.950 49.820 ;
        RECT 0.650 46.460 0.700 48.180 ;
        RECT 4.300 46.460 295.700 48.180 ;
        RECT 0.650 44.820 298.950 46.460 ;
        RECT 0.650 43.100 0.700 44.820 ;
        RECT 4.300 43.100 295.700 44.820 ;
        RECT 0.650 38.100 298.950 43.100 ;
        RECT 0.650 36.380 0.700 38.100 ;
        RECT 4.300 36.380 295.700 38.100 ;
        RECT 0.650 34.740 298.950 36.380 ;
        RECT 0.650 33.020 0.700 34.740 ;
        RECT 4.300 33.020 295.700 34.740 ;
        RECT 0.650 31.380 298.950 33.020 ;
        RECT 0.650 29.660 0.700 31.380 ;
        RECT 4.300 29.660 295.700 31.380 ;
        RECT 0.650 28.020 298.950 29.660 ;
        RECT 0.650 26.300 0.700 28.020 ;
        RECT 4.300 26.300 295.700 28.020 ;
        RECT 0.650 24.660 298.950 26.300 ;
        RECT 0.650 22.940 0.700 24.660 ;
        RECT 4.300 22.940 295.700 24.660 ;
        RECT 0.650 21.300 298.950 22.940 ;
        RECT 0.650 19.580 0.700 21.300 ;
        RECT 4.300 19.580 295.700 21.300 ;
        RECT 0.650 17.940 298.950 19.580 ;
        RECT 0.650 16.220 0.700 17.940 ;
        RECT 4.300 16.220 295.700 17.940 ;
        RECT 0.650 14.580 298.950 16.220 ;
        RECT 0.650 12.860 0.700 14.580 ;
        RECT 4.300 12.860 295.700 14.580 ;
        RECT 0.650 11.220 298.950 12.860 ;
        RECT 0.650 9.500 0.700 11.220 ;
        RECT 4.300 9.500 295.700 11.220 ;
        RECT 0.650 7.860 298.950 9.500 ;
        RECT 0.650 6.140 0.700 7.860 ;
        RECT 4.300 6.140 295.700 7.860 ;
        RECT 0.650 4.500 298.950 6.140 ;
        RECT 0.650 2.780 0.700 4.500 ;
        RECT 4.300 2.780 295.700 4.500 ;
        RECT 0.650 1.140 298.950 2.780 ;
        RECT 0.650 0.700 295.700 1.140 ;
      LAYER Metal4 ;
        RECT 263.900 243.130 264.180 252.470 ;
  END
END top_wrapper
END LIBRARY

